module SCM16 (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_Program # (.UUID(64'd3036675205634735936 ^ UUID), .WORD_WIDTH(64'd16), .DEFAULT_FILE_NAME("Program_2A247002B2183F40.w16.bin"), .ARG_SIG("Program_2A247002B2183F40=%s")) Program_0 (.clk(clk), .rst(rst), .address(wire_174), .out0(wire_26), .out1(wire_133), .out2(wire_112), .out3(wire_25));
  TC_Counter # (.UUID(64'd3613463651816973605 ^ UUID), .BIT_WIDTH(64'd16), .count(16'd4)) Counter16_1 (.clk(clk), .rst(rst), .save(wire_129), .in(wire_195), .out(wire_174));
  TC_Ram # (.UUID(64'd3779316721177258366 ^ UUID), .WORD_WIDTH(64'd16), .WORD_COUNT(64'd32768)) Ram_2 (.clk(clk), .rst(rst), .load(wire_77), .save(wire_191), .address({{16{1'b0}}, wire_45 }), .in0({{48{1'b0}}, wire_39 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_8_0), .out1(), .out2(), .out3());
  TC_Splitter16 # (.UUID(64'd1964885700083813915 ^ UUID)) Splitter16_3 (.in(wire_26[15:0]), .out0(), .out1(wire_181));
  TC_Splitter8 # (.UUID(64'd2865909427779811686 ^ UUID)) Splitter8_4 (.in(wire_183), .out0(), .out1(), .out2(), .out3(), .out4(wire_116), .out5(wire_190), .out6(wire_89), .out7(wire_66));
  TC_Register # (.UUID(64'd1768297580719965166 ^ UUID), .BIT_WIDTH(64'd16)) Register16_5 (.clk(clk), .rst(rst), .load(wire_230), .save(wire_147), .in(wire_8[15:0]), .out(wire_131));
  TC_Register # (.UUID(64'd12270441446668041 ^ UUID), .BIT_WIDTH(64'd16)) Register16_6 (.clk(clk), .rst(rst), .load(wire_186), .save(wire_70), .in(wire_8[15:0]), .out(wire_24));
  TC_Register # (.UUID(64'd3602252881066521773 ^ UUID), .BIT_WIDTH(64'd16)) Register16_7 (.clk(clk), .rst(rst), .load(wire_219), .save(wire_117), .in(wire_8[15:0]), .out(wire_98));
  TC_Register # (.UUID(64'd937036284257795972 ^ UUID), .BIT_WIDTH(64'd16)) Register16_8 (.clk(clk), .rst(rst), .load(wire_32), .save(wire_94), .in(wire_8[15:0]), .out(wire_86));
  TC_Register # (.UUID(64'd1771485704314964723 ^ UUID), .BIT_WIDTH(64'd16)) Register16_9 (.clk(clk), .rst(rst), .load(wire_88), .save(wire_177), .in(wire_8[15:0]), .out(wire_194));
  TC_Register # (.UUID(64'd1030977193978425972 ^ UUID), .BIT_WIDTH(64'd16)) Register16_10 (.clk(clk), .rst(rst), .load(wire_16), .save(wire_49), .in(wire_8[15:0]), .out(wire_7));
  TC_Register # (.UUID(64'd1897207591897939717 ^ UUID), .BIT_WIDTH(64'd16)) Register16_11 (.clk(clk), .rst(rst), .load(wire_175), .save(wire_136), .in(wire_8[15:0]), .out(wire_158));
  TC_Splitter16 # (.UUID(64'd1676756795661497062 ^ UUID)) Splitter16_12 (.in(wire_133[15:0]), .out0(wire_223), .out1());
  TC_Splitter16 # (.UUID(64'd2723123645093883319 ^ UUID)) Splitter16_13 (.in(wire_112[15:0]), .out0(wire_121), .out1());
  TC_Or # (.UUID(64'd3489109707031568152 ^ UUID), .BIT_WIDTH(64'd1)) Or_14 (.in0(wire_55), .in1(wire_140), .out(wire_166));
  TC_Or # (.UUID(64'd2757568662684548394 ^ UUID), .BIT_WIDTH(64'd1)) Or_15 (.in0(wire_99), .in1(wire_36), .out(wire_230));
  TC_Or # (.UUID(64'd2444150779797091056 ^ UUID), .BIT_WIDTH(64'd1)) Or_16 (.in0(wire_198), .in1(wire_0), .out(wire_186));
  TC_Or # (.UUID(64'd3998494940572441480 ^ UUID), .BIT_WIDTH(64'd1)) Or_17 (.in0(wire_18), .in1(wire_71), .out(wire_219));
  TC_Or # (.UUID(64'd3745487864523206918 ^ UUID), .BIT_WIDTH(64'd1)) Or_18 (.in0(wire_67), .in1(wire_78), .out(wire_32));
  TC_Or # (.UUID(64'd151306593792916243 ^ UUID), .BIT_WIDTH(64'd1)) Or_19 (.in0(wire_6), .in1(wire_170), .out(wire_88));
  TC_Or # (.UUID(64'd3493104666195700629 ^ UUID), .BIT_WIDTH(64'd1)) Or_20 (.in0(wire_59), .in1(wire_51), .out(wire_16));
  TC_Or # (.UUID(64'd3870924515638343503 ^ UUID), .BIT_WIDTH(64'd1)) Or_21 (.in0(wire_162), .in1(wire_42), .out(wire_175));
  TC_Splitter8 # (.UUID(64'd2466557324773763251 ^ UUID)) Splitter8_22 (.in(wire_223), .out0(wire_38), .out1(wire_148), .out2(wire_229), .out3(wire_224), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd1977466255751035882 ^ UUID)) Splitter8_23 (.in(wire_121), .out0(wire_153), .out1(wire_203), .out2(wire_105), .out3(wire_205), .out4(), .out5(), .out6(), .out7());
  TC_Splitter16 # (.UUID(64'd2261501443814513651 ^ UUID)) Splitter16_24 (.in(wire_25[15:0]), .out0(wire_215), .out1());
  TC_Splitter8 # (.UUID(64'd2576232014769382965 ^ UUID)) Splitter8_25 (.in(wire_215), .out0(wire_187), .out1(wire_168), .out2(wire_155), .out3(wire_179), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd2608661849516270155 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_26 (.en(wire_140), .in(wire_28), .out(wire_39_11));
  TC_Switch # (.UUID(64'd746143341221514145 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_27 (.en(wire_55), .in(wire_28), .out(wire_48_10));
  TC_Switch # (.UUID(64'd2038162143482139082 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_28 (.en(wire_36), .in(wire_131), .out(wire_39_10));
  TC_Switch # (.UUID(64'd4451929975376370007 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_29 (.en(wire_99), .in(wire_131), .out(wire_48_8));
  TC_Switch # (.UUID(64'd2149760867058136119 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_30 (.en(wire_0), .in(wire_24), .out(wire_39_9));
  TC_Switch # (.UUID(64'd1120920137235279511 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_31 (.en(wire_198), .in(wire_24), .out(wire_48_6));
  TC_Switch # (.UUID(64'd1049077220225763239 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_32 (.en(wire_71), .in(wire_98), .out(wire_39_8));
  TC_Switch # (.UUID(64'd690331529650965982 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_33 (.en(wire_18), .in(wire_98), .out(wire_48_4));
  TC_Switch # (.UUID(64'd4446234359163774586 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_34 (.en(wire_78), .in(wire_86), .out(wire_39_7));
  TC_Switch # (.UUID(64'd68561501764135042 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_35 (.en(wire_67), .in(wire_86), .out(wire_48_2));
  TC_Switch # (.UUID(64'd2300663947791505692 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_36 (.en(wire_170), .in(wire_194), .out(wire_39_6));
  TC_Switch # (.UUID(64'd1809390294038489791 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_37 (.en(wire_6), .in(wire_194), .out(wire_48_0));
  TC_Switch # (.UUID(64'd2131531128077507626 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_38 (.en(wire_51), .in(wire_7), .out(wire_39_5));
  TC_Switch # (.UUID(64'd2315389642693555300 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_39 (.en(wire_59), .in(wire_7), .out(wire_48_1));
  TC_Switch # (.UUID(64'd4187739606022409523 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_40 (.en(wire_42), .in(wire_158), .out(wire_39_4));
  TC_Switch # (.UUID(64'd1859071114078130426 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_41 (.en(wire_162), .in(wire_158), .out(wire_48_3));
  TC_Equal # (.UUID(64'd137163679941758477 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_42 (.in0(wire_26[15:0]), .in1(wire_202), .out(wire_74));
  TC_Halt # (.UUID(64'd2683931794444888664 ^ UUID)) Halt_43 (.clk(clk), .rst(rst), .en(wire_74));
  TC_Constant # (.UUID(64'd1352990490392554841 ^ UUID), .BIT_WIDTH(64'd16), .value(16'hFFFF)) Constant16_44 (.out(wire_202));
  TC_Switch # (.UUID(64'd971606683869478136 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_45 (.en(wire_89), .in(wire_112[15:0]), .out(wire_39_12));
  TC_Switch # (.UUID(64'd488700789590138722 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_46 (.en(wire_66), .in(wire_133[15:0]), .out(wire_48_12));
  TC_Constant # (.UUID(64'd1219804294531623130 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h0)) Constant16_47 (.out(wire_28));
  TC_Switch # (.UUID(64'd2854432665896608476 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_48 (.en(wire_50), .in(wire_181), .out(wire_183));
  TC_Not # (.UUID(64'd1919204710248089503 ^ UUID), .BIT_WIDTH(64'd1)) Not_49 (.in(wire_74), .out(wire_50));
  TC_Switch # (.UUID(64'd3648642341737646920 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_50 (.en(wire_129), .in(wire_25[15:0]), .out(wire_195));
  TC_Switch # (.UUID(64'd2839537485959427856 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_51 (.en(wire_97), .in(wire_97), .out(wire_129));
  TC_Splitter16 # (.UUID(64'd4451072885120255536 ^ UUID)) Splitter16_52 (.in(wire_26[15:0]), .out0(wire_208), .out1());
  TC_Splitter8 # (.UUID(64'd1191888651688547656 ^ UUID)) Splitter8_53 (.in(wire_208), .out0(wire_232), .out1(wire_200), .out2(wire_204), .out3(wire_111), .out4(), .out5(), .out6(), .out7());
  TC_Not # (.UUID(64'd4189336834672528069 ^ UUID), .BIT_WIDTH(64'd1)) Not_54 (.in(wire_63), .out(wire_138));
  TC_Add # (.UUID(64'd3182557287143411779 ^ UUID), .BIT_WIDTH(64'd16)) Add16_55 (.in0(wire_48), .in1(wire_39), .ci(1'd0), .out(wire_211), .co());
  TC_Add # (.UUID(64'd1424675120960351269 ^ UUID), .BIT_WIDTH(64'd16)) Add16_56 (.in0(wire_48), .in1(wire_25[15:0]), .ci(1'd0), .out(wire_80), .co());
  TC_Switch # (.UUID(64'd284020542177892273 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_57 (.en(wire_57), .in(wire_211), .out(wire_45_1));
  TC_Switch # (.UUID(64'd1034703434088870431 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_58 (.en(wire_125), .in(wire_80), .out(wire_45_0));
  TC_Or # (.UUID(64'd657814780105628035 ^ UUID), .BIT_WIDTH(64'd1)) Or_59 (.in0(wire_97), .in1(wire_125), .out(wire_213));
  TC_Console # (.UUID(64'd1550364046122691923 ^ UUID)) Console_60 (.clk(clk), .rst(rst), .offset({{16{1'b0}}, wire_84 }));
  TC_Ram # (.UUID(64'd2067412014399195219 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd65536)) Ram_61 (.clk(clk), .rst(rst), .load(1'd0), .save(wire_234), .address({{16{1'b0}}, wire_48 }), .in0({{48{1'b0}}, wire_39 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(), .out1(), .out2(), .out3());
  TC_Ram # (.UUID(64'd2804227458846121453 ^ UUID), .WORD_WIDTH(64'd16), .WORD_COUNT(64'd32768)) Ram_62 (.clk(clk), .rst(rst), .load(wire_134), .save(wire_45[0:0]), .address({{16{1'b0}}, wire_39 }), .in0(64'd0), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(), .out1(), .out2(), .out3());
  TC_Splitter16 # (.UUID(64'd763171029710359662 ^ UUID)) Splitter16_63 (.in(wire_45), .out0(), .out1(wire_206));
  TC_Splitter8 # (.UUID(64'd3824024877144842064 ^ UUID)) Splitter8_64 (.in(wire_206), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7(wire_152));
  TC_Decoder1 # (.UUID(64'd4576965811034017994 ^ UUID)) Decoder1_65 (.sel(wire_152), .out0(wire_9), .out1(wire_157));
  TC_Switch # (.UUID(64'd2746301141431459897 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_66 (.en(wire_9), .in(wire_125), .out(wire_191));
  TC_Switch # (.UUID(64'd3430101359472696647 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_67 (.en(wire_9), .in(wire_57), .out(wire_77));
  TC_Switch # (.UUID(64'd1728891745001622010 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_68 (.en(wire_157), .in(wire_57), .out(wire_182));
  TC_Switch # (.UUID(64'd4375680025586519226 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_69 (.en(wire_157), .in(wire_125), .out(wire_134));
  TC_Register # (.UUID(64'd2693553474459199961 ^ UUID), .BIT_WIDTH(64'd16)) Register16_70 (.clk(clk), .rst(rst), .load(wire_72), .save(wire_58), .in(wire_167), .out(wire_84));
  TC_Add # (.UUID(64'd3809269893433252203 ^ UUID), .BIT_WIDTH(64'd16)) Add16_71 (.in0(wire_84), .in1(wire_142), .ci(1'd0), .out(wire_167), .co());
  TC_Constant # (.UUID(64'd2151188605745524424 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_72 (.out(wire_72));
  TC_Constant # (.UUID(64'd1918094738540249611 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h50)) Constant16_73 (.out(wire_142));
  TC_Splitter16 # (.UUID(64'd4494426812884145071 ^ UUID)) Splitter16_74 (.in(wire_26[15:0]), .out0(wire_47), .out1());
  TC_Splitter8 # (.UUID(64'd1684985711211094078 ^ UUID)) Splitter8_75 (.in(wire_47), .out0(wire_143), .out1(wire_122), .out2(wire_172), .out3(wire_104), .out4(), .out5(), .out6(), .out7());
  TC_Not # (.UUID(64'd2891551810552540629 ^ UUID), .BIT_WIDTH(64'd1)) Not_76 (.in(wire_44), .out(wire_68));
  TC_Register # (.UUID(64'd3266843945445956355 ^ UUID), .BIT_WIDTH(64'd16)) Register16_77 (.clk(clk), .rst(rst), .load(wire_92), .save(wire_150), .in(wire_8[15:0]), .out(wire_108));
  TC_Register # (.UUID(64'd373441705232759894 ^ UUID), .BIT_WIDTH(64'd16)) Register16_78 (.clk(clk), .rst(rst), .load(wire_96), .save(wire_60), .in(wire_8[15:0]), .out(wire_226));
  TC_Register # (.UUID(64'd898762616312898673 ^ UUID), .BIT_WIDTH(64'd16)) Register16_79 (.clk(clk), .rst(rst), .load(wire_54), .save(wire_33), .in(wire_8[15:0]), .out(wire_188));
  TC_Register # (.UUID(64'd35259159018310512 ^ UUID), .BIT_WIDTH(64'd16)) Register16_80 (.clk(clk), .rst(rst), .load(wire_34), .save(wire_159), .in(wire_8[15:0]), .out(wire_192));
  TC_Or # (.UUID(64'd3408749404784824565 ^ UUID), .BIT_WIDTH(64'd1)) Or_81 (.in0(wire_64), .in1(wire_161), .out(wire_92));
  TC_Or # (.UUID(64'd2045434085000650231 ^ UUID), .BIT_WIDTH(64'd1)) Or_82 (.in0(wire_119), .in1(wire_103), .out(wire_96));
  TC_Or # (.UUID(64'd4235778316917593708 ^ UUID), .BIT_WIDTH(64'd1)) Or_83 (.in0(wire_81), .in1(wire_52), .out(wire_54));
  TC_Or # (.UUID(64'd1881922342948910945 ^ UUID), .BIT_WIDTH(64'd1)) Or_84 (.in0(wire_163), .in1(wire_61), .out(wire_34));
  TC_Switch # (.UUID(64'd3154836780073834162 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_85 (.en(wire_161), .in(wire_108), .out(wire_39_3));
  TC_Switch # (.UUID(64'd3206739131565530044 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_86 (.en(wire_64), .in(wire_108), .out(wire_48_5));
  TC_Switch # (.UUID(64'd1476550871400967823 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_87 (.en(wire_103), .in(wire_226), .out(wire_39_2));
  TC_Switch # (.UUID(64'd1622071797847061869 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_88 (.en(wire_119), .in(wire_226), .out(wire_48_7));
  TC_Switch # (.UUID(64'd189967047438908968 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_89 (.en(wire_52), .in(wire_188), .out(wire_39_1));
  TC_Switch # (.UUID(64'd3142169352616083849 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_90 (.en(wire_81), .in(wire_188), .out(wire_48_9));
  TC_Switch # (.UUID(64'd2790449206563351533 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_91 (.en(wire_61), .in(wire_192), .out(wire_39_0));
  TC_Switch # (.UUID(64'd1382504743536358321 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_92 (.en(wire_163), .in(wire_192), .out(wire_48_11));
  TC_DotMatrixDisplay # (.UUID(64'd2660535027850879501 ^ UUID)) DotMatrixDisplay_93 (.clk(clk), .rst(rst), .en_y(wire_46[0:0]), .en_x(wire_20[0:0]), .color_info(wire_46[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd1287415170352733091 ^ UUID)) DotMatrixDisplay_94 (.clk(clk), .rst(rst), .en_y(wire_79[0:0]), .en_x(wire_20[0:0]), .color_info(wire_79[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd4375632836552484410 ^ UUID)) DotMatrixDisplay_95 (.clk(clk), .rst(rst), .en_y(wire_91[0:0]), .en_x(wire_20[0:0]), .color_info(wire_91[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd4352128498737539568 ^ UUID)) DotMatrixDisplay_96 (.clk(clk), .rst(rst), .en_y(wire_93[0:0]), .en_x(wire_20[0:0]), .color_info(wire_93[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd4375805759909017124 ^ UUID)) DotMatrixDisplay_97 (.clk(clk), .rst(rst), .en_y(wire_5[0:0]), .en_x(wire_20[0:0]), .color_info(wire_5[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd4001708814053949966 ^ UUID)) DotMatrixDisplay_98 (.clk(clk), .rst(rst), .en_y(wire_30[0:0]), .en_x(wire_20[0:0]), .color_info(wire_30[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd3789421783879759989 ^ UUID)) DotMatrixDisplay_99 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_20[0:0]), .color_info(wire_23[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd3949917514357280402 ^ UUID)) DotMatrixDisplay_100 (.clk(clk), .rst(rst), .en_y(wire_29[0:0]), .en_x(wire_3[0:0]), .color_info(wire_29[31:0]), .pixel_info(wire_3));
  TC_DotMatrixDisplay # (.UUID(64'd1120366264718111392 ^ UUID)) DotMatrixDisplay_101 (.clk(clk), .rst(rst), .en_y(wire_46[0:0]), .en_x(wire_3[0:0]), .color_info(wire_46[31:0]), .pixel_info(wire_3));
  TC_DotMatrixDisplay # (.UUID(64'd3830190475406040627 ^ UUID)) DotMatrixDisplay_102 (.clk(clk), .rst(rst), .en_y(wire_79[0:0]), .en_x(wire_3[0:0]), .color_info(wire_79[31:0]), .pixel_info(wire_3));
  TC_DotMatrixDisplay # (.UUID(64'd3695649649918959220 ^ UUID)) DotMatrixDisplay_103 (.clk(clk), .rst(rst), .en_y(wire_91[0:0]), .en_x(wire_3[0:0]), .color_info(wire_91[31:0]), .pixel_info(wire_3));
  TC_DotMatrixDisplay # (.UUID(64'd2190167902128485018 ^ UUID)) DotMatrixDisplay_104 (.clk(clk), .rst(rst), .en_y(wire_93[0:0]), .en_x(wire_3[0:0]), .color_info(wire_93[31:0]), .pixel_info(wire_3));
  TC_DotMatrixDisplay # (.UUID(64'd108023444932811778 ^ UUID)) DotMatrixDisplay_105 (.clk(clk), .rst(rst), .en_y(wire_93[0:0]), .en_x(wire_2[0:0]), .color_info(wire_93[31:0]), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd3127548314519555293 ^ UUID)) DotMatrixDisplay_106 (.clk(clk), .rst(rst), .en_y(wire_5[0:0]), .en_x(wire_3[0:0]), .color_info(wire_5[31:0]), .pixel_info(wire_3));
  TC_DotMatrixDisplay # (.UUID(64'd3232957164641830670 ^ UUID)) DotMatrixDisplay_107 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_3[0:0]), .color_info(wire_23[31:0]), .pixel_info(wire_3));
  TC_DotMatrixDisplay # (.UUID(64'd2013870924499775536 ^ UUID)) DotMatrixDisplay_108 (.clk(clk), .rst(rst), .en_y(wire_29[0:0]), .en_x(wire_2[0:0]), .color_info(wire_29[31:0]), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd1700230642759998846 ^ UUID)) DotMatrixDisplay_109 (.clk(clk), .rst(rst), .en_y(wire_46[0:0]), .en_x(wire_2[0:0]), .color_info(wire_46[31:0]), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd640862205653523348 ^ UUID)) DotMatrixDisplay_110 (.clk(clk), .rst(rst), .en_y(wire_79[0:0]), .en_x(wire_2[0:0]), .color_info(wire_79[31:0]), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd1441056504049384023 ^ UUID)) DotMatrixDisplay_111 (.clk(clk), .rst(rst), .en_y(wire_91[0:0]), .en_x(wire_2[0:0]), .color_info(wire_91[31:0]), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd4360991051994526462 ^ UUID)) DotMatrixDisplay_112 (.clk(clk), .rst(rst), .en_y(wire_93[0:0]), .en_x(wire_35[0:0]), .color_info(wire_93[31:0]), .pixel_info(wire_35));
  TC_DotMatrixDisplay # (.UUID(64'd3732720467344721449 ^ UUID)) DotMatrixDisplay_113 (.clk(clk), .rst(rst), .en_y(wire_30[0:0]), .en_x(wire_3[0:0]), .color_info(wire_30[31:0]), .pixel_info(wire_3));
  TC_DotMatrixDisplay # (.UUID(64'd3164120181411694497 ^ UUID)) DotMatrixDisplay_114 (.clk(clk), .rst(rst), .en_y(wire_30[0:0]), .en_x(wire_2[0:0]), .color_info(wire_30[31:0]), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd3058994005473620099 ^ UUID)) DotMatrixDisplay_115 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_2[0:0]), .color_info(wire_23[31:0]), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd3043865689462340485 ^ UUID)) DotMatrixDisplay_116 (.clk(clk), .rst(rst), .en_y(wire_29[0:0]), .en_x(wire_35[0:0]), .color_info(wire_29[31:0]), .pixel_info(wire_35));
  TC_DotMatrixDisplay # (.UUID(64'd1232256408208860842 ^ UUID)) DotMatrixDisplay_117 (.clk(clk), .rst(rst), .en_y(wire_46[0:0]), .en_x(wire_35[0:0]), .color_info(wire_46[31:0]), .pixel_info(wire_35));
  TC_DotMatrixDisplay # (.UUID(64'd456775015865694566 ^ UUID)) DotMatrixDisplay_118 (.clk(clk), .rst(rst), .en_y(wire_79[0:0]), .en_x(wire_35[0:0]), .color_info(wire_79[31:0]), .pixel_info(wire_35));
  TC_DotMatrixDisplay # (.UUID(64'd1486947349792475943 ^ UUID)) DotMatrixDisplay_119 (.clk(clk), .rst(rst), .en_y(wire_91[0:0]), .en_x(wire_35[0:0]), .color_info(wire_91[31:0]), .pixel_info(wire_35));
  TC_DotMatrixDisplay # (.UUID(64'd1986390658814520529 ^ UUID)) DotMatrixDisplay_120 (.clk(clk), .rst(rst), .en_y(wire_5[0:0]), .en_x(wire_2[0:0]), .color_info(wire_5[31:0]), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd428599916565265934 ^ UUID)) DotMatrixDisplay_121 (.clk(clk), .rst(rst), .en_y(wire_5[0:0]), .en_x(wire_35[0:0]), .color_info(wire_5[31:0]), .pixel_info(wire_35));
  TC_DotMatrixDisplay # (.UUID(64'd1361741769374930265 ^ UUID)) DotMatrixDisplay_122 (.clk(clk), .rst(rst), .en_y(wire_30[0:0]), .en_x(wire_35[0:0]), .color_info(wire_30[31:0]), .pixel_info(wire_35));
  TC_DotMatrixDisplay # (.UUID(64'd3810902491231665649 ^ UUID)) DotMatrixDisplay_123 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_35[0:0]), .color_info(wire_23[31:0]), .pixel_info(wire_35));
  TC_DotMatrixDisplay # (.UUID(64'd145789043302394905 ^ UUID)) DotMatrixDisplay_124 (.clk(clk), .rst(rst), .en_y(wire_29[0:0]), .en_x(wire_19[0:0]), .color_info(wire_29[31:0]), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd3780736919653097053 ^ UUID)) DotMatrixDisplay_125 (.clk(clk), .rst(rst), .en_y(wire_46[0:0]), .en_x(wire_19[0:0]), .color_info(wire_46[31:0]), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd2485800408185936591 ^ UUID)) DotMatrixDisplay_126 (.clk(clk), .rst(rst), .en_y(wire_79[0:0]), .en_x(wire_19[0:0]), .color_info(wire_79[31:0]), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd3637982062020866444 ^ UUID)) DotMatrixDisplay_127 (.clk(clk), .rst(rst), .en_y(wire_91[0:0]), .en_x(wire_19[0:0]), .color_info(wire_91[31:0]), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd2077992963286351604 ^ UUID)) DotMatrixDisplay_128 (.clk(clk), .rst(rst), .en_y(wire_93[0:0]), .en_x(wire_19[0:0]), .color_info(wire_93[31:0]), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd3780255053339576859 ^ UUID)) DotMatrixDisplay_129 (.clk(clk), .rst(rst), .en_y(wire_5[0:0]), .en_x(wire_19[0:0]), .color_info(wire_5[31:0]), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd3088612785393467744 ^ UUID)) DotMatrixDisplay_130 (.clk(clk), .rst(rst), .en_y(wire_30[0:0]), .en_x(wire_19[0:0]), .color_info(wire_30[31:0]), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd4340287621202113208 ^ UUID)) DotMatrixDisplay_131 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_19[0:0]), .color_info(wire_23[31:0]), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd3263142337545802511 ^ UUID)) DotMatrixDisplay_132 (.clk(clk), .rst(rst), .en_y(wire_29[0:0]), .en_x(wire_1[0:0]), .color_info(wire_29[31:0]), .pixel_info(wire_1));
  TC_DotMatrixDisplay # (.UUID(64'd4368304585025255821 ^ UUID)) DotMatrixDisplay_133 (.clk(clk), .rst(rst), .en_y(wire_46[0:0]), .en_x(wire_1[0:0]), .color_info(wire_46[31:0]), .pixel_info(wire_1));
  TC_DotMatrixDisplay # (.UUID(64'd3035154864325599620 ^ UUID)) DotMatrixDisplay_134 (.clk(clk), .rst(rst), .en_y(wire_79[0:0]), .en_x(wire_1[0:0]), .color_info(wire_79[31:0]), .pixel_info(wire_1));
  TC_DotMatrixDisplay # (.UUID(64'd1984067145119237049 ^ UUID)) DotMatrixDisplay_135 (.clk(clk), .rst(rst), .en_y(wire_91[0:0]), .en_x(wire_1[0:0]), .color_info(wire_91[31:0]), .pixel_info(wire_1));
  TC_DotMatrixDisplay # (.UUID(64'd257903097512365689 ^ UUID)) DotMatrixDisplay_136 (.clk(clk), .rst(rst), .en_y(wire_93[0:0]), .en_x(wire_1[0:0]), .color_info(wire_93[31:0]), .pixel_info(wire_1));
  TC_DotMatrixDisplay # (.UUID(64'd1855803350615582069 ^ UUID)) DotMatrixDisplay_137 (.clk(clk), .rst(rst), .en_y(wire_5[0:0]), .en_x(wire_1[0:0]), .color_info(wire_5[31:0]), .pixel_info(wire_1));
  TC_DotMatrixDisplay # (.UUID(64'd4156190447566119276 ^ UUID)) DotMatrixDisplay_138 (.clk(clk), .rst(rst), .en_y(wire_30[0:0]), .en_x(wire_1[0:0]), .color_info(wire_30[31:0]), .pixel_info(wire_1));
  TC_DotMatrixDisplay # (.UUID(64'd3549196530068966916 ^ UUID)) DotMatrixDisplay_139 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_1[0:0]), .color_info(wire_23[31:0]), .pixel_info(wire_1));
  TC_SegmentDisplay # (.UUID(64'd4189100092568263645 ^ UUID)) SegmentDisplay_140 (.clk(clk), .rst(rst), .enable(wire_56), .value(8'd0));
  TC_SegmentDisplay # (.UUID(64'd736833738424528830 ^ UUID)) SegmentDisplay_141 (.clk(clk), .rst(rst), .enable(wire_56), .value(8'd0));
  TC_SegmentDisplay # (.UUID(64'd2349681992692057466 ^ UUID)) SegmentDisplay_142 (.clk(clk), .rst(rst), .enable(wire_56), .value(8'd0));
  TC_SegmentDisplay # (.UUID(64'd3433535943137751453 ^ UUID)) SegmentDisplay_143 (.clk(clk), .rst(rst), .enable(wire_56), .value(8'd0));
  TC_SegmentDisplay # (.UUID(64'd3098309455346325270 ^ UUID)) SegmentDisplay_144 (.clk(clk), .rst(rst), .enable(wire_56), .value(8'd0));
  TC_Constant # (.UUID(64'd430758642605415045 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_145 (.out(wire_56));
  TC_DotMatrixDisplay # (.UUID(64'd3746276803240527606 ^ UUID)) DotMatrixDisplay_146 (.clk(clk), .rst(rst), .en_y(wire_29[0:0]), .en_x(wire_20[0:0]), .color_info(wire_29[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd4237472817339994162 ^ UUID)) DotMatrixDisplay_147 (.clk(clk), .rst(rst), .en_y(wire_37[0:0]), .en_x(wire_20[0:0]), .color_info(wire_37[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd1177830180225486220 ^ UUID)) DotMatrixDisplay_148 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_20[0:0]), .color_info(wire_73[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd250680188831281298 ^ UUID)) DotMatrixDisplay_149 (.clk(clk), .rst(rst), .en_y(wire_41[0:0]), .en_x(wire_20[0:0]), .color_info(wire_41[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd1576462328986410349 ^ UUID)) DotMatrixDisplay_150 (.clk(clk), .rst(rst), .en_y(wire_10[0:0]), .en_x(wire_20[0:0]), .color_info(wire_10[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd316625153349409673 ^ UUID)) DotMatrixDisplay_151 (.clk(clk), .rst(rst), .en_y(wire_11[0:0]), .en_x(wire_20[0:0]), .color_info(wire_11[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd959143668139620378 ^ UUID)) DotMatrixDisplay_152 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_20[0:0]), .color_info(wire_13[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd684938010714015909 ^ UUID)) DotMatrixDisplay_153 (.clk(clk), .rst(rst), .en_y(wire_126[0:0]), .en_x(wire_20[0:0]), .color_info(wire_126[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd1796769576252909689 ^ UUID)) DotMatrixDisplay_154 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_3[0:0]), .color_info(wire_40[31:0]), .pixel_info(wire_3));
  TC_DotMatrixDisplay # (.UUID(64'd28266181691657389 ^ UUID)) DotMatrixDisplay_155 (.clk(clk), .rst(rst), .en_y(wire_37[0:0]), .en_x(wire_3[0:0]), .color_info(wire_37[31:0]), .pixel_info(wire_3));
  TC_DotMatrixDisplay # (.UUID(64'd3196962412568546329 ^ UUID)) DotMatrixDisplay_156 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_3[0:0]), .color_info(wire_73[31:0]), .pixel_info(wire_3));
  TC_DotMatrixDisplay # (.UUID(64'd2205871638966640606 ^ UUID)) DotMatrixDisplay_157 (.clk(clk), .rst(rst), .en_y(wire_41[0:0]), .en_x(wire_3[0:0]), .color_info(wire_41[31:0]), .pixel_info(wire_3));
  TC_DotMatrixDisplay # (.UUID(64'd3874186372446959361 ^ UUID)) DotMatrixDisplay_158 (.clk(clk), .rst(rst), .en_y(wire_10[0:0]), .en_x(wire_3[0:0]), .color_info(wire_10[31:0]), .pixel_info(wire_3));
  TC_DotMatrixDisplay # (.UUID(64'd2720360903878823189 ^ UUID)) DotMatrixDisplay_159 (.clk(clk), .rst(rst), .en_y(wire_11[0:0]), .en_x(wire_3[0:0]), .color_info(wire_11[31:0]), .pixel_info(wire_3));
  TC_DotMatrixDisplay # (.UUID(64'd504346027738870704 ^ UUID)) DotMatrixDisplay_160 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_3[0:0]), .color_info(wire_13[31:0]), .pixel_info(wire_3));
  TC_DotMatrixDisplay # (.UUID(64'd184655924988308158 ^ UUID)) DotMatrixDisplay_161 (.clk(clk), .rst(rst), .en_y(wire_126[0:0]), .en_x(wire_3[0:0]), .color_info(wire_126[31:0]), .pixel_info(wire_3));
  TC_DotMatrixDisplay # (.UUID(64'd3162126675592577790 ^ UUID)) DotMatrixDisplay_162 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_2[0:0]), .color_info(wire_40[31:0]), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd841957664227372441 ^ UUID)) DotMatrixDisplay_163 (.clk(clk), .rst(rst), .en_y(wire_37[0:0]), .en_x(wire_2[0:0]), .color_info(wire_37[31:0]), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd4388146087367304388 ^ UUID)) DotMatrixDisplay_164 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_2[0:0]), .color_info(wire_73[31:0]), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd935756330229132165 ^ UUID)) DotMatrixDisplay_165 (.clk(clk), .rst(rst), .en_y(wire_41[0:0]), .en_x(wire_2[0:0]), .color_info(wire_41[31:0]), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd38018604794773973 ^ UUID)) DotMatrixDisplay_166 (.clk(clk), .rst(rst), .en_y(wire_10[0:0]), .en_x(wire_2[0:0]), .color_info(wire_10[31:0]), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd1334297701942639290 ^ UUID)) DotMatrixDisplay_167 (.clk(clk), .rst(rst), .en_y(wire_11[0:0]), .en_x(wire_2[0:0]), .color_info(wire_11[31:0]), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd971239419644370685 ^ UUID)) DotMatrixDisplay_168 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_2[0:0]), .color_info(wire_13[31:0]), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd2299276613863097833 ^ UUID)) DotMatrixDisplay_169 (.clk(clk), .rst(rst), .en_y(wire_126[0:0]), .en_x(wire_2[0:0]), .color_info(wire_126[31:0]), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd4066308585007913895 ^ UUID)) DotMatrixDisplay_170 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_35[0:0]), .color_info(wire_40[31:0]), .pixel_info(wire_35));
  TC_DotMatrixDisplay # (.UUID(64'd1188730429928185190 ^ UUID)) DotMatrixDisplay_171 (.clk(clk), .rst(rst), .en_y(wire_37[0:0]), .en_x(wire_35[0:0]), .color_info(wire_37[31:0]), .pixel_info(wire_35));
  TC_DotMatrixDisplay # (.UUID(64'd4280800355417676313 ^ UUID)) DotMatrixDisplay_172 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_35[0:0]), .color_info(wire_73[31:0]), .pixel_info(wire_35));
  TC_DotMatrixDisplay # (.UUID(64'd4360520332522264149 ^ UUID)) DotMatrixDisplay_173 (.clk(clk), .rst(rst), .en_y(wire_41[0:0]), .en_x(wire_35[0:0]), .color_info(wire_41[31:0]), .pixel_info(wire_35));
  TC_DotMatrixDisplay # (.UUID(64'd475575386071264203 ^ UUID)) DotMatrixDisplay_174 (.clk(clk), .rst(rst), .en_y(wire_10[0:0]), .en_x(wire_35[0:0]), .color_info(wire_10[31:0]), .pixel_info(wire_35));
  TC_DotMatrixDisplay # (.UUID(64'd4099921249160036118 ^ UUID)) DotMatrixDisplay_175 (.clk(clk), .rst(rst), .en_y(wire_11[0:0]), .en_x(wire_35[0:0]), .color_info(wire_11[31:0]), .pixel_info(wire_35));
  TC_DotMatrixDisplay # (.UUID(64'd2008157871612466016 ^ UUID)) DotMatrixDisplay_176 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_35[0:0]), .color_info(wire_13[31:0]), .pixel_info(wire_35));
  TC_DotMatrixDisplay # (.UUID(64'd3526081255155773975 ^ UUID)) DotMatrixDisplay_177 (.clk(clk), .rst(rst), .en_y(wire_126[0:0]), .en_x(wire_35[0:0]), .color_info(wire_126[31:0]), .pixel_info(wire_35));
  TC_DotMatrixDisplay # (.UUID(64'd1085763782026657154 ^ UUID)) DotMatrixDisplay_178 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_19[0:0]), .color_info(wire_40[31:0]), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd1935004646604641077 ^ UUID)) DotMatrixDisplay_179 (.clk(clk), .rst(rst), .en_y(wire_37[0:0]), .en_x(wire_19[0:0]), .color_info(wire_37[31:0]), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd4228153944513970773 ^ UUID)) DotMatrixDisplay_180 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_19[0:0]), .color_info(wire_73[31:0]), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd3380853135653261586 ^ UUID)) DotMatrixDisplay_181 (.clk(clk), .rst(rst), .en_y(wire_41[0:0]), .en_x(wire_19[0:0]), .color_info(wire_41[31:0]), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd142464094186867413 ^ UUID)) DotMatrixDisplay_182 (.clk(clk), .rst(rst), .en_y(wire_10[0:0]), .en_x(wire_19[0:0]), .color_info(wire_10[31:0]), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd988217888803392985 ^ UUID)) DotMatrixDisplay_183 (.clk(clk), .rst(rst), .en_y(wire_11[0:0]), .en_x(wire_19[0:0]), .color_info(wire_11[31:0]), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd54720530278277779 ^ UUID)) DotMatrixDisplay_184 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_19[0:0]), .color_info(wire_13[31:0]), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd2688678971804628028 ^ UUID)) DotMatrixDisplay_185 (.clk(clk), .rst(rst), .en_y(wire_126[0:0]), .en_x(wire_19[0:0]), .color_info(wire_126[31:0]), .pixel_info(wire_19));
  TC_DotMatrixDisplay # (.UUID(64'd553058778145918310 ^ UUID)) DotMatrixDisplay_186 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_1[0:0]), .color_info(wire_40[31:0]), .pixel_info(wire_1));
  TC_DotMatrixDisplay # (.UUID(64'd2098597773896322169 ^ UUID)) DotMatrixDisplay_187 (.clk(clk), .rst(rst), .en_y(wire_37[0:0]), .en_x(wire_1[0:0]), .color_info(wire_37[31:0]), .pixel_info(wire_1));
  TC_DotMatrixDisplay # (.UUID(64'd1919740307961683958 ^ UUID)) DotMatrixDisplay_188 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_1[0:0]), .color_info(wire_73[31:0]), .pixel_info(wire_1));
  TC_DotMatrixDisplay # (.UUID(64'd2955390637246533656 ^ UUID)) DotMatrixDisplay_189 (.clk(clk), .rst(rst), .en_y(wire_41[0:0]), .en_x(wire_1[0:0]), .color_info(wire_41[31:0]), .pixel_info(wire_1));
  TC_DotMatrixDisplay # (.UUID(64'd3399628396733223633 ^ UUID)) DotMatrixDisplay_190 (.clk(clk), .rst(rst), .en_y(wire_10[0:0]), .en_x(wire_1[0:0]), .color_info(wire_10[31:0]), .pixel_info(wire_1));
  TC_DotMatrixDisplay # (.UUID(64'd1503255611657110166 ^ UUID)) DotMatrixDisplay_191 (.clk(clk), .rst(rst), .en_y(wire_11[0:0]), .en_x(wire_1[0:0]), .color_info(wire_11[31:0]), .pixel_info(wire_1));
  TC_DotMatrixDisplay # (.UUID(64'd1934210770642016723 ^ UUID)) DotMatrixDisplay_192 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_1[0:0]), .color_info(wire_13[31:0]), .pixel_info(wire_1));
  TC_DotMatrixDisplay # (.UUID(64'd4430890296674284431 ^ UUID)) DotMatrixDisplay_193 (.clk(clk), .rst(rst), .en_y(wire_126[0:0]), .en_x(wire_1[0:0]), .color_info(wire_126[31:0]), .pixel_info(wire_1));
  TC_DotMatrixDisplay # (.UUID(64'd1370192036403734636 ^ UUID)) DotMatrixDisplay_194 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_20[0:0]), .color_info(wire_40[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd1914293527285665104 ^ UUID)) DotMatrixDisplay_195 (.clk(clk), .rst(rst), .en_y(wire_29[0:0]), .en_x(wire_17[0:0]), .color_info(wire_29[31:0]), .pixel_info(wire_17));
  TC_DotMatrixDisplay # (.UUID(64'd4024378624965788820 ^ UUID)) DotMatrixDisplay_196 (.clk(clk), .rst(rst), .en_y(wire_46[0:0]), .en_x(wire_17[0:0]), .color_info(wire_46[31:0]), .pixel_info(wire_17));
  TC_DotMatrixDisplay # (.UUID(64'd331796838499445221 ^ UUID)) DotMatrixDisplay_197 (.clk(clk), .rst(rst), .en_y(wire_79[0:0]), .en_x(wire_17[0:0]), .color_info(wire_79[31:0]), .pixel_info(wire_17));
  TC_DotMatrixDisplay # (.UUID(64'd1109146203016946320 ^ UUID)) DotMatrixDisplay_198 (.clk(clk), .rst(rst), .en_y(wire_91[0:0]), .en_x(wire_17[0:0]), .color_info(wire_91[31:0]), .pixel_info(wire_17));
  TC_DotMatrixDisplay # (.UUID(64'd2037862037394616530 ^ UUID)) DotMatrixDisplay_199 (.clk(clk), .rst(rst), .en_y(wire_93[0:0]), .en_x(wire_17[0:0]), .color_info(wire_93[31:0]), .pixel_info(wire_17));
  TC_DotMatrixDisplay # (.UUID(64'd756317346051932726 ^ UUID)) DotMatrixDisplay_200 (.clk(clk), .rst(rst), .en_y(wire_5[0:0]), .en_x(wire_17[0:0]), .color_info(wire_5[31:0]), .pixel_info(wire_17));
  TC_DotMatrixDisplay # (.UUID(64'd741221856880638315 ^ UUID)) DotMatrixDisplay_201 (.clk(clk), .rst(rst), .en_y(wire_30[0:0]), .en_x(wire_17[0:0]), .color_info(wire_30[31:0]), .pixel_info(wire_17));
  TC_DotMatrixDisplay # (.UUID(64'd2554897745454830451 ^ UUID)) DotMatrixDisplay_202 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_17[0:0]), .color_info(wire_23[31:0]), .pixel_info(wire_17));
  TC_DotMatrixDisplay # (.UUID(64'd4352234980297914729 ^ UUID)) DotMatrixDisplay_203 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_17[0:0]), .color_info(wire_40[31:0]), .pixel_info(wire_17));
  TC_DotMatrixDisplay # (.UUID(64'd4044674900922762564 ^ UUID)) DotMatrixDisplay_204 (.clk(clk), .rst(rst), .en_y(wire_37[0:0]), .en_x(wire_17[0:0]), .color_info(wire_37[31:0]), .pixel_info(wire_17));
  TC_DotMatrixDisplay # (.UUID(64'd2175572511635428388 ^ UUID)) DotMatrixDisplay_205 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_17[0:0]), .color_info(wire_73[31:0]), .pixel_info(wire_17));
  TC_DotMatrixDisplay # (.UUID(64'd1352766524066348872 ^ UUID)) DotMatrixDisplay_206 (.clk(clk), .rst(rst), .en_y(wire_41[0:0]), .en_x(wire_17[0:0]), .color_info(wire_41[31:0]), .pixel_info(wire_17));
  TC_DotMatrixDisplay # (.UUID(64'd1625039672493008527 ^ UUID)) DotMatrixDisplay_207 (.clk(clk), .rst(rst), .en_y(wire_10[0:0]), .en_x(wire_17[0:0]), .color_info(wire_10[31:0]), .pixel_info(wire_17));
  TC_DotMatrixDisplay # (.UUID(64'd672361543425103183 ^ UUID)) DotMatrixDisplay_208 (.clk(clk), .rst(rst), .en_y(wire_11[0:0]), .en_x(wire_17[0:0]), .color_info(wire_11[31:0]), .pixel_info(wire_17));
  TC_DotMatrixDisplay # (.UUID(64'd1607234245481583786 ^ UUID)) DotMatrixDisplay_209 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_17[0:0]), .color_info(wire_13[31:0]), .pixel_info(wire_17));
  TC_DotMatrixDisplay # (.UUID(64'd2377050978244241774 ^ UUID)) DotMatrixDisplay_210 (.clk(clk), .rst(rst), .en_y(wire_126[0:0]), .en_x(wire_17[0:0]), .color_info(wire_126[31:0]), .pixel_info(wire_17));
  TC_DotMatrixDisplay # (.UUID(64'd3222873545553085433 ^ UUID)) DotMatrixDisplay_211 (.clk(clk), .rst(rst), .en_y(wire_29[0:0]), .en_x(wire_4[0:0]), .color_info(wire_29[31:0]), .pixel_info(wire_4));
  TC_DotMatrixDisplay # (.UUID(64'd3188765738163086443 ^ UUID)) DotMatrixDisplay_212 (.clk(clk), .rst(rst), .en_y(wire_46[0:0]), .en_x(wire_4[0:0]), .color_info(wire_46[31:0]), .pixel_info(wire_4));
  TC_DotMatrixDisplay # (.UUID(64'd838700140978907233 ^ UUID)) DotMatrixDisplay_213 (.clk(clk), .rst(rst), .en_y(wire_79[0:0]), .en_x(wire_4[0:0]), .color_info(wire_79[31:0]), .pixel_info(wire_4));
  TC_DotMatrixDisplay # (.UUID(64'd3920730297055212015 ^ UUID)) DotMatrixDisplay_214 (.clk(clk), .rst(rst), .en_y(wire_91[0:0]), .en_x(wire_4[0:0]), .color_info(wire_91[31:0]), .pixel_info(wire_4));
  TC_DotMatrixDisplay # (.UUID(64'd3481948759443637 ^ UUID)) DotMatrixDisplay_215 (.clk(clk), .rst(rst), .en_y(wire_93[0:0]), .en_x(wire_4[0:0]), .color_info(wire_93[31:0]), .pixel_info(wire_4));
  TC_DotMatrixDisplay # (.UUID(64'd511172518486640794 ^ UUID)) DotMatrixDisplay_216 (.clk(clk), .rst(rst), .en_y(wire_5[0:0]), .en_x(wire_4[0:0]), .color_info(wire_5[31:0]), .pixel_info(wire_4));
  TC_DotMatrixDisplay # (.UUID(64'd4053020964562097569 ^ UUID)) DotMatrixDisplay_217 (.clk(clk), .rst(rst), .en_y(wire_30[0:0]), .en_x(wire_4[0:0]), .color_info(wire_30[31:0]), .pixel_info(wire_4));
  TC_DotMatrixDisplay # (.UUID(64'd3303805443456392646 ^ UUID)) DotMatrixDisplay_218 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_4[0:0]), .color_info(wire_23[31:0]), .pixel_info(wire_4));
  TC_DotMatrixDisplay # (.UUID(64'd3229541704842781328 ^ UUID)) DotMatrixDisplay_219 (.clk(clk), .rst(rst), .en_y(wire_40[0:0]), .en_x(wire_4[0:0]), .color_info(wire_40[31:0]), .pixel_info(wire_4));
  TC_DotMatrixDisplay # (.UUID(64'd1520258463232062736 ^ UUID)) DotMatrixDisplay_220 (.clk(clk), .rst(rst), .en_y(wire_37[0:0]), .en_x(wire_4[0:0]), .color_info(wire_37[31:0]), .pixel_info(wire_4));
  TC_DotMatrixDisplay # (.UUID(64'd3535073739167951615 ^ UUID)) DotMatrixDisplay_221 (.clk(clk), .rst(rst), .en_y(wire_73[0:0]), .en_x(wire_4[0:0]), .color_info(wire_73[31:0]), .pixel_info(wire_4));
  TC_DotMatrixDisplay # (.UUID(64'd2508590195121546232 ^ UUID)) DotMatrixDisplay_222 (.clk(clk), .rst(rst), .en_y(wire_41[0:0]), .en_x(wire_4[0:0]), .color_info(wire_41[31:0]), .pixel_info(wire_4));
  TC_DotMatrixDisplay # (.UUID(64'd4190156087276806644 ^ UUID)) DotMatrixDisplay_223 (.clk(clk), .rst(rst), .en_y(wire_10[0:0]), .en_x(wire_4[0:0]), .color_info(wire_10[31:0]), .pixel_info(wire_4));
  TC_DotMatrixDisplay # (.UUID(64'd3357160141127693591 ^ UUID)) DotMatrixDisplay_224 (.clk(clk), .rst(rst), .en_y(wire_11[0:0]), .en_x(wire_4[0:0]), .color_info(wire_11[31:0]), .pixel_info(wire_4));
  TC_DotMatrixDisplay # (.UUID(64'd3712829154125709738 ^ UUID)) DotMatrixDisplay_225 (.clk(clk), .rst(rst), .en_y(wire_13[0:0]), .en_x(wire_4[0:0]), .color_info(wire_13[31:0]), .pixel_info(wire_4));
  TC_DotMatrixDisplay # (.UUID(64'd2545725033216246256 ^ UUID)) DotMatrixDisplay_226 (.clk(clk), .rst(rst), .en_y(wire_126[0:0]), .en_x(wire_4[0:0]), .color_info(wire_126[31:0]), .pixel_info(wire_4));
  TC_Mul # (.UUID(64'd2748524405844472327 ^ UUID), .BIT_WIDTH(64'd16)) DivMod16_227 (.in0(wire_39), .in1(wire_214), .out0(wire_100), .out1(wire_114));
  TC_Mul # (.UUID(64'd4020347048163863131 ^ UUID), .BIT_WIDTH(64'd16)) DivMod16_228 (.in0(wire_48), .in1(wire_235), .out0(wire_173), .out1(wire_62));
  TC_Constant # (.UUID(64'd1313141643564538265 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h6)) Constant16_229 (.out(wire_235));
  TC_Constant # (.UUID(64'd4112089032370153264 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h8)) Constant16_230 (.out(wire_214));
  TC_Splitter16 # (.UUID(64'd2668786745693159507 ^ UUID)) Splitter16_231 (.in(wire_173), .out0(wire_184), .out1());
  TC_Splitter8 # (.UUID(64'd2631886754935636255 ^ UUID)) Splitter8_232 (.in(wire_184), .out0(wire_217), .out1(wire_218), .out2(wire_43), .out3(wire_83), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd550414518326034956 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_233 (.en(wire_165), .in(wire_12), .out(wire_29));
  TC_Switch # (.UUID(64'd977382900955430648 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_234 (.en(wire_176), .in(wire_12), .out(wire_46));
  TC_Switch # (.UUID(64'd1891242292111482311 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_235 (.en(wire_149), .in(wire_12), .out(wire_79));
  TC_Switch # (.UUID(64'd856889246029500943 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_236 (.en(wire_27), .in(wire_12), .out(wire_91));
  TC_Switch # (.UUID(64'd3189954206832060770 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_237 (.en(wire_127), .in(wire_12), .out(wire_93));
  TC_Switch # (.UUID(64'd2600416908798528202 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_238 (.en(wire_90), .in(wire_12), .out(wire_5));
  TC_Switch # (.UUID(64'd3352059561228947819 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_239 (.en(wire_123), .in(wire_12), .out(wire_30));
  TC_Switch # (.UUID(64'd3576546926653500711 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_240 (.en(wire_87), .in(wire_12), .out(wire_23));
  TC_Switch # (.UUID(64'd773945265408688934 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_241 (.en(wire_15), .in(wire_12), .out(wire_40));
  TC_Switch # (.UUID(64'd4124677947420211807 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_242 (.en(wire_130), .in(wire_12), .out(wire_37));
  TC_Switch # (.UUID(64'd1892597805610563739 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_243 (.en(wire_135), .in(wire_12), .out(wire_73));
  TC_Switch # (.UUID(64'd4501036839557111240 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_244 (.en(wire_22), .in(wire_12), .out(wire_41));
  TC_Switch # (.UUID(64'd2653282250793028984 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_245 (.en(wire_110), .in(wire_12), .out(wire_10));
  TC_Switch # (.UUID(64'd2835551167096927095 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_246 (.en(wire_151), .in(wire_12), .out(wire_11));
  TC_Switch # (.UUID(64'd811538821685340963 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_247 (.en(wire_76), .in(wire_12), .out(wire_13));
  TC_Switch # (.UUID(64'd1795419328706358879 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_248 (.en(wire_132), .in(wire_12), .out(wire_126));
  TC_Switch # (.UUID(64'd3384031002647223712 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_249 (.en(wire_85), .in(wire_75), .out(wire_20));
  TC_Switch # (.UUID(64'd796360369331162321 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_250 (.en(wire_107), .in(wire_75), .out(wire_3));
  TC_Switch # (.UUID(64'd770893388854325356 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_251 (.en(wire_139), .in(wire_75), .out(wire_2));
  TC_Switch # (.UUID(64'd2296729005521048932 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_252 (.en(wire_180), .in(wire_75), .out(wire_35));
  TC_Switch # (.UUID(64'd2700874401252926434 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_253 (.en(wire_109), .in(wire_75), .out(wire_19));
  TC_Switch # (.UUID(64'd3871697537247032043 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_254 (.en(wire_193), .in(wire_75), .out(wire_1));
  TC_Switch # (.UUID(64'd1657382633537052929 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_255 (.en(wire_209), .in(wire_75), .out(wire_17));
  TC_Switch # (.UUID(64'd2430440528996199989 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_256 (.en(wire_82), .in(wire_75), .out(wire_4));
  TC_Mul # (.UUID(64'd1323562681874756164 ^ UUID), .BIT_WIDTH(64'd16)) Mul16_257 (.in0(wire_114), .in1(wire_221), .out0(wire_197), .out1());
  TC_Constant # (.UUID(64'd625362193213988375 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h6)) Constant16_258 (.out(wire_221));
  TC_Add # (.UUID(64'd4099861895360639395 ^ UUID), .BIT_WIDTH(64'd16)) Add16_259 (.in0(wire_62), .in1(wire_65), .ci(1'd0), .out(wire_101), .co());
  TC_Constant # (.UUID(64'd3900858799247905575 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h8)) Constant16_260 (.out(wire_216));
  TC_Constant # (.UUID(64'd2454158573449235377 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h1)) Constant16_261 (.out(wire_212));
  TC_Shl # (.UUID(64'd191663886776180221 ^ UUID), .BIT_WIDTH(64'd64)) Shl64_262 (.in({{48{1'b0}}, wire_212 }), .shift(wire_101[7:0]), .out(wire_171));
  TC_Or # (.UUID(64'd3463268789363960265 ^ UUID), .BIT_WIDTH(64'd64)) Or64_263 (.in0(wire_171), .in1(wire_141), .out(wire_222));
  TC_Constant # (.UUID(64'd213891297043897909 ^ UUID), .BIT_WIDTH(64'd64), .value(64'h100000000000001)) Constant64_264 (.out(wire_141));
  TC_Splitter8 # (.UUID(64'd4038412651713004570 ^ UUID)) Splitter8_265 (.in(wire_233), .out0(wire_160), .out1(wire_201), .out2(wire_21), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter16 # (.UUID(64'd3776431078096079195 ^ UUID)) Splitter16_266 (.in(wire_100), .out0(wire_233), .out1());
  TC_Decoder3 # (.UUID(64'd4013734321313478962 ^ UUID)) Decoder3_267 (.dis(1'd0), .sel0(wire_160), .sel1(wire_201), .sel2(wire_21), .out0(wire_220), .out1(wire_169), .out2(wire_137), .out3(wire_102), .out4(wire_146), .out5(wire_53), .out6(wire_144), .out7(wire_128));
  TC_Maker64 # (.UUID(64'd1192448886920089561 ^ UUID)) Maker64_268 (.in0(wire_227), .in1(wire_145), .in2(wire_225), .in3(wire_178), .in4(8'd0), .in5(8'd0), .in6(8'd0), .in7(8'd0), .out(wire_12));
  TC_Constant # (.UUID(64'd803552191146308597 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h34)) Constant8_269 (.out(wire_178));
  TC_Constant # (.UUID(64'd511943185350590578 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h77)) Constant8_270 (.out(wire_225));
  TC_Constant # (.UUID(64'd222105970335437196 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hEB)) Constant8_271 (.out(wire_145));
  TC_Add # (.UUID(64'd2037122097572093298 ^ UUID), .BIT_WIDTH(64'd16)) Add16_272 (.in0(wire_197), .in1(wire_216), .ci(1'd0), .out(wire_65), .co());
  DEC4 # (.UUID(64'd606098422439323267 ^ UUID)) DEC4_273 (.clk(clk), .rst(rst), .Bit_1(wire_38), .Bit_2(wire_148), .Bit_3(wire_229), .Bit_4(wire_224), .Disable(wire_66), .Output_1(wire_6), .Output_2(wire_59), .Output_3(wire_162), .Output_4(wire_67), .Output_5(wire_18), .Output_6(wire_198), .Output_7(wire_99), .Output_8(wire_55), .Output_9(wire_64), .Output_10(wire_119), .Output_11(wire_81), .Output_12(wire_163), .Output_13(), .Output_14(), .Output_15(), .Output_16());
  DEC4 # (.UUID(64'd2350125178974466839 ^ UUID)) DEC4_274 (.clk(clk), .rst(rst), .Bit_1(wire_153), .Bit_2(wire_203), .Bit_3(wire_105), .Bit_4(wire_205), .Disable(wire_89), .Output_1(wire_170), .Output_2(wire_51), .Output_3(wire_42), .Output_4(wire_78), .Output_5(wire_71), .Output_6(wire_0), .Output_7(wire_36), .Output_8(wire_140), .Output_9(wire_161), .Output_10(wire_103), .Output_11(wire_52), .Output_12(wire_61), .Output_13(), .Output_14(), .Output_15(), .Output_16());
  DEC4 # (.UUID(64'd4239434022177334522 ^ UUID)) DEC4_275 (.clk(clk), .rst(rst), .Bit_1(wire_187), .Bit_2(wire_168), .Bit_3(wire_155), .Bit_4(wire_179), .Disable(wire_213), .Output_1(wire_177), .Output_2(wire_49), .Output_3(wire_136), .Output_4(wire_94), .Output_5(wire_117), .Output_6(wire_70), .Output_7(wire_147), .Output_8(wire_156), .Output_9(wire_150), .Output_10(wire_60), .Output_11(wire_33), .Output_12(wire_159), .Output_13(), .Output_14(), .Output_15(), .Output_16());
  DEC2 # (.UUID(64'd2289023201248810830 ^ UUID)) DEC2_276 (.clk(clk), .rst(rst), .Input_1(wire_116), .Input_2(wire_190), .Disable(wire_74), .Output_1(wire_95), .Output_2(wire_63), .Output_3(wire_44), .Output_4(wire_31));
  DEC4 # (.UUID(64'd2197146422829533631 ^ UUID)) DEC4_277 (.clk(clk), .rst(rst), .Bit_1(wire_232), .Bit_2(wire_200), .Bit_3(wire_204), .Bit_4(wire_111), .Disable(wire_138), .Output_1(), .Output_2(), .Output_3(), .Output_4(), .Output_5(), .Output_6(), .Output_7(wire_125), .Output_8(wire_57), .Output_9(), .Output_10(), .Output_11(), .Output_12(), .Output_13(), .Output_14(), .Output_15(), .Output_16());
  ALU # (.UUID(64'd2893949216972807263 ^ UUID)) ALU_278 (.clk(clk), .rst(rst), .Instruction(wire_26[15:0]), .Input_1(wire_48), .Input_2(wire_39), .Enable(wire_31), .Output(wire_8_1[15:0]));
  COND # (.UUID(64'd1476889620975298455 ^ UUID)) COND_279 (.clk(clk), .rst(rst), .Instruction(wire_26[15:0]), .Input_1(wire_48), .Input_2(wire_39), .Enable(wire_95), .Output(wire_97));
  DEC4 # (.UUID(64'd2773479126471196673 ^ UUID)) DEC4_280 (.clk(clk), .rst(rst), .Bit_1(wire_143), .Bit_2(wire_122), .Bit_3(wire_172), .Bit_4(wire_104), .Disable(wire_68), .Output_1(), .Output_2(), .Output_3(), .Output_4(), .Output_5(wire_164), .Output_6(wire_124), .Output_7(wire_58), .Output_8(wire_234), .Output_9(), .Output_10(), .Output_11(), .Output_12(), .Output_13(), .Output_14(), .Output_15(), .Output_16());
  DEC4 # (.UUID(64'd302757758434011087 ^ UUID)) DEC4_281 (.clk(clk), .rst(rst), .Bit_1(wire_217), .Bit_2(wire_218), .Bit_3(wire_43), .Bit_4(wire_83), .Disable(1'd0), .Output_1(wire_207), .Output_2(wire_196), .Output_3(wire_228), .Output_4(wire_113), .Output_5(wire_106), .Output_6(wire_210), .Output_7(wire_185), .Output_8(wire_69), .Output_9(wire_14), .Output_10(wire_231), .Output_11(wire_120), .Output_12(wire_199), .Output_13(wire_189), .Output_14(wire_154), .Output_15(wire_118), .Output_16(wire_115));
  OPP16 # (.UUID(64'd319281544511355177 ^ UUID)) OPP16_282 (.clk(clk), .rst(rst), .Input_1(wire_69), .Input_2(wire_185), .Input_3(wire_210), .Input_4(wire_106), .Input_5(wire_113), .Input_6(wire_207), .Input_7(wire_196), .Input_8(wire_228), .Input_9(wire_14), .Input_10(wire_231), .Input_11(wire_120), .Input_12(wire_199), .Input_13(wire_189), .Input_14(wire_154), .Input_15(wire_118), .Input_16(wire_115), .Output_1(wire_132), .Output_2(wire_76), .Output_3(wire_151), .Output_4(wire_110), .Output_5(wire_22), .Output_6(wire_135), .Output_7(wire_130), .Output_8(wire_15), .Output_9(wire_87), .Output_10(wire_123), .Output_11(wire_90), .Output_12(wire_127), .Output_13(wire_27), .Output_14(wire_149), .Output_15(wire_176), .Output_16(wire_165));
  OPP8 # (.UUID(64'd3315969898736290245 ^ UUID)) OPP8_283 (.clk(clk), .rst(rst), .Input_1(wire_220), .Input_2(wire_169), .Input_3(wire_137), .Input_4(wire_102), .Input_5(wire_146), .Input_6(wire_53), .Input_7(wire_144), .Input_8(wire_128), .Output_1(wire_85), .Output_2(wire_107), .Output_3(wire_139), .Output_4(wire_180), .Output_5(wire_109), .Output_6(wire_193), .Output_7(wire_209), .Output_8(wire_82));
  TC_Mux # (.UUID(64'd3182122184138242733 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_284 (.sel(wire_124), .in0(64'd0), .in1(wire_222), .out(wire_75));
  TC_Constant # (.UUID(64'd499839709284412840 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_285 (.out(wire_227));

  wire [0:0] wire_0;
  wire [63:0] wire_1;
  wire [63:0] wire_2;
  wire [63:0] wire_3;
  wire [63:0] wire_4;
  wire [63:0] wire_5;
  wire [0:0] wire_6;
  wire [15:0] wire_7;
  wire [63:0] wire_8;
  wire [63:0] wire_8_0;
  wire [63:0] wire_8_1;
  assign wire_8 = wire_8_0|wire_8_1;
  wire [0:0] wire_9;
  wire [63:0] wire_10;
  wire [63:0] wire_11;
  wire [63:0] wire_12;
  wire [63:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [63:0] wire_17;
  wire [0:0] wire_18;
  wire [63:0] wire_19;
  wire [63:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [63:0] wire_23;
  wire [15:0] wire_24;
  wire [63:0] wire_25;
  wire [63:0] wire_26;
  wire [0:0] wire_27;
  wire [15:0] wire_28;
  wire [63:0] wire_29;
  wire [63:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [63:0] wire_35;
  wire [0:0] wire_36;
  wire [63:0] wire_37;
  wire [0:0] wire_38;
  wire [15:0] wire_39;
  wire [15:0] wire_39_0;
  wire [15:0] wire_39_1;
  wire [15:0] wire_39_2;
  wire [15:0] wire_39_3;
  wire [15:0] wire_39_4;
  wire [15:0] wire_39_5;
  wire [15:0] wire_39_6;
  wire [15:0] wire_39_7;
  wire [15:0] wire_39_8;
  wire [15:0] wire_39_9;
  wire [15:0] wire_39_10;
  wire [15:0] wire_39_11;
  wire [15:0] wire_39_12;
  assign wire_39 = wire_39_0|wire_39_1|wire_39_2|wire_39_3|wire_39_4|wire_39_5|wire_39_6|wire_39_7|wire_39_8|wire_39_9|wire_39_10|wire_39_11|wire_39_12;
  wire [63:0] wire_40;
  wire [63:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;
  wire [15:0] wire_45;
  wire [15:0] wire_45_0;
  wire [15:0] wire_45_1;
  assign wire_45 = wire_45_0|wire_45_1;
  wire [63:0] wire_46;
  wire [7:0] wire_47;
  wire [15:0] wire_48;
  wire [15:0] wire_48_0;
  wire [15:0] wire_48_1;
  wire [15:0] wire_48_2;
  wire [15:0] wire_48_3;
  wire [15:0] wire_48_4;
  wire [15:0] wire_48_5;
  wire [15:0] wire_48_6;
  wire [15:0] wire_48_7;
  wire [15:0] wire_48_8;
  wire [15:0] wire_48_9;
  wire [15:0] wire_48_10;
  wire [15:0] wire_48_11;
  wire [15:0] wire_48_12;
  assign wire_48 = wire_48_0|wire_48_1|wire_48_2|wire_48_3|wire_48_4|wire_48_5|wire_48_6|wire_48_7|wire_48_8|wire_48_9|wire_48_10|wire_48_11|wire_48_12;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [0:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [15:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  wire [15:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [0:0] wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [63:0] wire_73;
  wire [0:0] wire_74;
  wire [63:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [63:0] wire_79;
  wire [15:0] wire_80;
  wire [0:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;
  wire [15:0] wire_84;
  wire [0:0] wire_85;
  wire [15:0] wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;
  wire [0:0] wire_90;
  wire [63:0] wire_91;
  wire [0:0] wire_92;
  wire [63:0] wire_93;
  wire [0:0] wire_94;
  wire [0:0] wire_95;
  wire [0:0] wire_96;
  wire [0:0] wire_97;
  wire [15:0] wire_98;
  wire [0:0] wire_99;
  wire [15:0] wire_100;
  wire [15:0] wire_101;
  wire [0:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [0:0] wire_105;
  wire [0:0] wire_106;
  wire [0:0] wire_107;
  wire [15:0] wire_108;
  wire [0:0] wire_109;
  wire [0:0] wire_110;
  wire [0:0] wire_111;
  wire [63:0] wire_112;
  wire [0:0] wire_113;
  wire [15:0] wire_114;
  wire [0:0] wire_115;
  wire [0:0] wire_116;
  wire [0:0] wire_117;
  wire [0:0] wire_118;
  wire [0:0] wire_119;
  wire [0:0] wire_120;
  wire [7:0] wire_121;
  wire [0:0] wire_122;
  wire [0:0] wire_123;
  wire [0:0] wire_124;
  wire [0:0] wire_125;
  wire [63:0] wire_126;
  wire [0:0] wire_127;
  wire [0:0] wire_128;
  wire [0:0] wire_129;
  wire [0:0] wire_130;
  wire [15:0] wire_131;
  wire [0:0] wire_132;
  wire [63:0] wire_133;
  wire [0:0] wire_134;
  wire [0:0] wire_135;
  wire [0:0] wire_136;
  wire [0:0] wire_137;
  wire [0:0] wire_138;
  wire [0:0] wire_139;
  wire [0:0] wire_140;
  wire [63:0] wire_141;
  wire [15:0] wire_142;
  wire [0:0] wire_143;
  wire [0:0] wire_144;
  wire [7:0] wire_145;
  wire [0:0] wire_146;
  wire [0:0] wire_147;
  wire [0:0] wire_148;
  wire [0:0] wire_149;
  wire [0:0] wire_150;
  wire [0:0] wire_151;
  wire [0:0] wire_152;
  wire [0:0] wire_153;
  wire [0:0] wire_154;
  wire [0:0] wire_155;
  wire [0:0] wire_156;
  wire [0:0] wire_157;
  wire [15:0] wire_158;
  wire [0:0] wire_159;
  wire [0:0] wire_160;
  wire [0:0] wire_161;
  wire [0:0] wire_162;
  wire [0:0] wire_163;
  wire [0:0] wire_164;
  wire [0:0] wire_165;
  wire [0:0] wire_166;
  wire [15:0] wire_167;
  wire [0:0] wire_168;
  wire [0:0] wire_169;
  wire [0:0] wire_170;
  wire [63:0] wire_171;
  wire [0:0] wire_172;
  wire [15:0] wire_173;
  wire [15:0] wire_174;
  wire [0:0] wire_175;
  wire [0:0] wire_176;
  wire [0:0] wire_177;
  wire [7:0] wire_178;
  wire [0:0] wire_179;
  wire [0:0] wire_180;
  wire [7:0] wire_181;
  wire [0:0] wire_182;
  wire [7:0] wire_183;
  wire [7:0] wire_184;
  wire [0:0] wire_185;
  wire [0:0] wire_186;
  wire [0:0] wire_187;
  wire [15:0] wire_188;
  wire [0:0] wire_189;
  wire [0:0] wire_190;
  wire [0:0] wire_191;
  wire [15:0] wire_192;
  wire [0:0] wire_193;
  wire [15:0] wire_194;
  wire [15:0] wire_195;
  wire [0:0] wire_196;
  wire [15:0] wire_197;
  wire [0:0] wire_198;
  wire [0:0] wire_199;
  wire [0:0] wire_200;
  wire [0:0] wire_201;
  wire [15:0] wire_202;
  wire [0:0] wire_203;
  wire [0:0] wire_204;
  wire [0:0] wire_205;
  wire [7:0] wire_206;
  wire [0:0] wire_207;
  wire [7:0] wire_208;
  wire [0:0] wire_209;
  wire [0:0] wire_210;
  wire [15:0] wire_211;
  wire [15:0] wire_212;
  wire [0:0] wire_213;
  wire [15:0] wire_214;
  wire [7:0] wire_215;
  wire [15:0] wire_216;
  wire [0:0] wire_217;
  wire [0:0] wire_218;
  wire [0:0] wire_219;
  wire [0:0] wire_220;
  wire [15:0] wire_221;
  wire [63:0] wire_222;
  wire [7:0] wire_223;
  wire [0:0] wire_224;
  wire [7:0] wire_225;
  wire [15:0] wire_226;
  wire [7:0] wire_227;
  wire [0:0] wire_228;
  wire [0:0] wire_229;
  wire [0:0] wire_230;
  wire [0:0] wire_231;
  wire [0:0] wire_232;
  wire [7:0] wire_233;
  wire [0:0] wire_234;
  wire [15:0] wire_235;

endmodule
