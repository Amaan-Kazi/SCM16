module OPP16 (clk, rst, Input_1, Input_2, Input_3, Input_4, Input_5, Input_6, Input_7, Input_8, Input_9, Input_10, Input_11, Input_12, Input_13, Input_14, Input_15, Input_16, Enable_All, Output_1, Output_2, Output_3, Output_4, Output_5, Output_6, Output_7, Output_8, Output_9, Output_10, Output_11, Output_12, Output_13, Output_14, Output_15, Output_16);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] Input_1;
  input  wire [0:0] Input_2;
  input  wire [0:0] Input_3;
  input  wire [0:0] Input_4;
  input  wire [0:0] Input_5;
  input  wire [0:0] Input_6;
  input  wire [0:0] Input_7;
  input  wire [0:0] Input_8;
  input  wire [0:0] Input_9;
  input  wire [0:0] Input_10;
  input  wire [0:0] Input_11;
  input  wire [0:0] Input_12;
  input  wire [0:0] Input_13;
  input  wire [0:0] Input_14;
  input  wire [0:0] Input_15;
  input  wire [0:0] Input_16;
  input  wire [0:0] Enable_All;
  output  wire [0:0] Output_1;
  output  wire [0:0] Output_2;
  output  wire [0:0] Output_3;
  output  wire [0:0] Output_4;
  output  wire [0:0] Output_5;
  output  wire [0:0] Output_6;
  output  wire [0:0] Output_7;
  output  wire [0:0] Output_8;
  output  wire [0:0] Output_9;
  output  wire [0:0] Output_10;
  output  wire [0:0] Output_11;
  output  wire [0:0] Output_12;
  output  wire [0:0] Output_13;
  output  wire [0:0] Output_14;
  output  wire [0:0] Output_15;
  output  wire [0:0] Output_16;

  TC_Maker16 # (.UUID(64'd4576894713119714030 ^ UUID)) Maker16_0 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd4159457257671284809 ^ UUID)) Maker16_1 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd135754618811469109 ^ UUID)) Maker16_2 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd2144888840407442937 ^ UUID)) Maker16_3 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd925366045232949744 ^ UUID)) Maker16_4 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd753355972069108851 ^ UUID)) Maker16_5 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd1697733420865645326 ^ UUID)) Maker16_6 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd923918180205380539 ^ UUID)) Maker16_7 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd3574614010472517973 ^ UUID)) Maker16_8 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd88510775329053771 ^ UUID)) Maker16_9 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd3562464275485822968 ^ UUID)) Maker16_10 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd2946293184664622310 ^ UUID)) Maker16_11 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd1923742623033063111 ^ UUID)) Maker16_12 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd2531585302615411283 ^ UUID)) Maker16_13 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd1446271324425451477 ^ UUID)) Maker16_14 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd971499438910037494 ^ UUID)) Maker16_15 (.in0(8'd0), .in1(8'd0), .out());
  TC_Or # (.UUID(64'd464374234935265593 ^ UUID), .BIT_WIDTH(64'd1)) Or_16 (.in0(wire_1), .in1(wire_0), .out(wire_14));
  TC_Or # (.UUID(64'd1487585136896219486 ^ UUID), .BIT_WIDTH(64'd1)) Or_17 (.in0(wire_1), .in1(wire_19), .out(wire_26));
  TC_Or # (.UUID(64'd129943381723371862 ^ UUID), .BIT_WIDTH(64'd1)) Or_18 (.in0(wire_1), .in1(wire_22), .out(wire_31));
  TC_Or # (.UUID(64'd1435292707242546051 ^ UUID), .BIT_WIDTH(64'd1)) Or_19 (.in0(wire_1), .in1(wire_6), .out(wire_11));
  TC_Or # (.UUID(64'd2403491923322782475 ^ UUID), .BIT_WIDTH(64'd1)) Or_20 (.in0(wire_1), .in1(wire_7), .out(wire_21));
  TC_Or # (.UUID(64'd2607232073358608135 ^ UUID), .BIT_WIDTH(64'd1)) Or_21 (.in0(wire_1), .in1(wire_18), .out(wire_28));
  TC_Or # (.UUID(64'd2764809654089472988 ^ UUID), .BIT_WIDTH(64'd1)) Or_22 (.in0(wire_1), .in1(wire_2), .out(wire_4));
  TC_Or # (.UUID(64'd2056166774136696565 ^ UUID), .BIT_WIDTH(64'd1)) Or_23 (.in0(wire_1), .in1(wire_9), .out(wire_27));
  TC_Or # (.UUID(64'd4539864918566049744 ^ UUID), .BIT_WIDTH(64'd1)) Or_24 (.in0(wire_1), .in1(wire_5), .out(wire_32));
  TC_Or # (.UUID(64'd4294436867348702187 ^ UUID), .BIT_WIDTH(64'd1)) Or_25 (.in0(wire_1), .in1(wire_16), .out(wire_8));
  TC_Or # (.UUID(64'd2651740742167582059 ^ UUID), .BIT_WIDTH(64'd1)) Or_26 (.in0(wire_1), .in1(wire_20), .out(wire_15));
  TC_Or # (.UUID(64'd1101571698995348906 ^ UUID), .BIT_WIDTH(64'd1)) Or_27 (.in0(wire_1), .in1(wire_17), .out(wire_24));
  TC_Or # (.UUID(64'd4575843383047068471 ^ UUID), .BIT_WIDTH(64'd1)) Or_28 (.in0(wire_1), .in1(wire_3), .out(wire_29));
  TC_Or # (.UUID(64'd3876158841287781865 ^ UUID), .BIT_WIDTH(64'd1)) Or_29 (.in0(wire_1), .in1(wire_25), .out(wire_23));
  TC_Or # (.UUID(64'd1988900315667371397 ^ UUID), .BIT_WIDTH(64'd1)) Or_30 (.in0(wire_1), .in1(wire_10), .out(wire_30));
  TC_Or # (.UUID(64'd4259045747919882354 ^ UUID), .BIT_WIDTH(64'd1)) Or_31 (.in0(wire_1), .in1(wire_12), .out(wire_13));

  wire [0:0] wire_0;
  assign wire_0 = Input_16;
  wire [0:0] wire_1;
  assign wire_1 = Enable_All;
  wire [0:0] wire_2;
  assign wire_2 = Input_10;
  wire [0:0] wire_3;
  assign wire_3 = Input_4;
  wire [0:0] wire_4;
  assign Output_7 = wire_4;
  wire [0:0] wire_5;
  assign wire_5 = Input_8;
  wire [0:0] wire_6;
  assign wire_6 = Input_13;
  wire [0:0] wire_7;
  assign wire_7 = Input_12;
  wire [0:0] wire_8;
  assign Output_10 = wire_8;
  wire [0:0] wire_9;
  assign wire_9 = Input_9;
  wire [0:0] wire_10;
  assign wire_10 = Input_2;
  wire [0:0] wire_11;
  assign Output_4 = wire_11;
  wire [0:0] wire_12;
  assign wire_12 = Input_1;
  wire [0:0] wire_13;
  assign Output_16 = wire_13;
  wire [0:0] wire_14;
  assign Output_1 = wire_14;
  wire [0:0] wire_15;
  assign Output_11 = wire_15;
  wire [0:0] wire_16;
  assign wire_16 = Input_7;
  wire [0:0] wire_17;
  assign wire_17 = Input_5;
  wire [0:0] wire_18;
  assign wire_18 = Input_11;
  wire [0:0] wire_19;
  assign wire_19 = Input_15;
  wire [0:0] wire_20;
  assign wire_20 = Input_6;
  wire [0:0] wire_21;
  assign Output_5 = wire_21;
  wire [0:0] wire_22;
  assign wire_22 = Input_14;
  wire [0:0] wire_23;
  assign Output_14 = wire_23;
  wire [0:0] wire_24;
  assign Output_12 = wire_24;
  wire [0:0] wire_25;
  assign wire_25 = Input_3;
  wire [0:0] wire_26;
  assign Output_2 = wire_26;
  wire [0:0] wire_27;
  assign Output_8 = wire_27;
  wire [0:0] wire_28;
  assign Output_6 = wire_28;
  wire [0:0] wire_29;
  assign Output_13 = wire_29;
  wire [0:0] wire_30;
  assign Output_15 = wire_30;
  wire [0:0] wire_31;
  assign Output_3 = wire_31;
  wire [0:0] wire_32;
  assign Output_9 = wire_32;

endmodule
