module SCM16 (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_Program # (.UUID(64'd3036675205634735936 ^ UUID), .WORD_WIDTH(64'd16), .DEFAULT_FILE_NAME("Program_2A247002B2183F40.w16.bin"), .ARG_SIG("Program_2A247002B2183F40=%s")) Program_0 (.clk(clk), .rst(rst), .address(wire_126), .out0(wire_97), .out1(wire_13), .out2(wire_95), .out3(wire_25));
  TC_Counter # (.UUID(64'd3613463651816973605 ^ UUID), .BIT_WIDTH(64'd16), .count(16'd4)) Counter16_1 (.clk(clk), .rst(rst), .save(wire_83), .in(wire_115), .out(wire_126));
  TC_Ram # (.UUID(64'd3779316721177258366 ^ UUID), .WORD_WIDTH(64'd16), .WORD_COUNT(64'd32768)) Ram_2 (.clk(clk), .rst(rst), .load(wire_170), .save(wire_235), .address({{16{1'b0}}, wire_93 }), .in0({{48{1'b0}}, wire_44 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_26_0), .out1(), .out2(), .out3());
  TC_Splitter16 # (.UUID(64'd1964885700083813915 ^ UUID)) Splitter16_3 (.in(wire_97[15:0]), .out0(), .out1(wire_189));
  TC_Splitter8 # (.UUID(64'd2865909427779811686 ^ UUID)) Splitter8_4 (.in(wire_260), .out0(), .out1(), .out2(), .out3(), .out4(wire_240), .out5(wire_176), .out6(wire_103), .out7(wire_124));
  TC_Register # (.UUID(64'd1768297580719965166 ^ UUID), .BIT_WIDTH(64'd16)) Register16_5 (.clk(clk), .rst(rst), .load(wire_173), .save(wire_150), .in(wire_26[15:0]), .out(wire_141));
  TC_Register # (.UUID(64'd12270441446668041 ^ UUID), .BIT_WIDTH(64'd16)) Register16_6 (.clk(clk), .rst(rst), .load(wire_163), .save(wire_205), .in(wire_26[15:0]), .out(wire_33));
  TC_Register # (.UUID(64'd3602252881066521773 ^ UUID), .BIT_WIDTH(64'd16)) Register16_7 (.clk(clk), .rst(rst), .load(wire_230), .save(wire_70), .in(wire_26[15:0]), .out(wire_147));
  TC_Register # (.UUID(64'd937036284257795972 ^ UUID), .BIT_WIDTH(64'd16)) Register16_8 (.clk(clk), .rst(rst), .load(wire_120), .save(wire_136), .in(wire_26[15:0]), .out(wire_161));
  TC_Register # (.UUID(64'd1771485704314964723 ^ UUID), .BIT_WIDTH(64'd16)) Register16_9 (.clk(clk), .rst(rst), .load(wire_245), .save(wire_73), .in(wire_26[15:0]), .out(wire_86));
  TC_Register # (.UUID(64'd1030977193978425972 ^ UUID), .BIT_WIDTH(64'd16)) Register16_10 (.clk(clk), .rst(rst), .load(wire_279), .save(wire_34), .in(wire_26[15:0]), .out(wire_138));
  TC_Register # (.UUID(64'd1897207591897939717 ^ UUID), .BIT_WIDTH(64'd16)) Register16_11 (.clk(clk), .rst(rst), .load(wire_128), .save(wire_74), .in(wire_26[15:0]), .out(wire_214));
  TC_Splitter16 # (.UUID(64'd1676756795661497062 ^ UUID)) Splitter16_12 (.in(wire_13[15:0]), .out0(wire_157), .out1());
  TC_Splitter16 # (.UUID(64'd2723123645093883319 ^ UUID)) Splitter16_13 (.in(wire_95[15:0]), .out0(wire_191), .out1());
  TC_Or # (.UUID(64'd3489109707031568152 ^ UUID), .BIT_WIDTH(64'd1)) Or_14 (.in0(wire_18), .in1(wire_50), .out(wire_265));
  TC_Or # (.UUID(64'd2757568662684548394 ^ UUID), .BIT_WIDTH(64'd1)) Or_15 (.in0(wire_8), .in1(wire_75), .out(wire_173));
  TC_Or # (.UUID(64'd2444150779797091056 ^ UUID), .BIT_WIDTH(64'd1)) Or_16 (.in0(wire_88), .in1(wire_106), .out(wire_163));
  TC_Or # (.UUID(64'd3998494940572441480 ^ UUID), .BIT_WIDTH(64'd1)) Or_17 (.in0(wire_139), .in1(wire_36), .out(wire_230));
  TC_Or # (.UUID(64'd3745487864523206918 ^ UUID), .BIT_WIDTH(64'd1)) Or_18 (.in0(wire_61), .in1(wire_179), .out(wire_120));
  TC_Or # (.UUID(64'd151306593792916243 ^ UUID), .BIT_WIDTH(64'd1)) Or_19 (.in0(wire_142), .in1(wire_38), .out(wire_245));
  TC_Or # (.UUID(64'd3493104666195700629 ^ UUID), .BIT_WIDTH(64'd1)) Or_20 (.in0(wire_42), .in1(wire_165), .out(wire_279));
  TC_Or # (.UUID(64'd3870924515638343503 ^ UUID), .BIT_WIDTH(64'd1)) Or_21 (.in0(wire_111), .in1(wire_114), .out(wire_128));
  TC_Splitter8 # (.UUID(64'd2466557324773763251 ^ UUID)) Splitter8_22 (.in(wire_157), .out0(wire_130), .out1(wire_185), .out2(wire_239), .out3(wire_277), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd1977466255751035882 ^ UUID)) Splitter8_23 (.in(wire_191), .out0(wire_216), .out1(wire_98), .out2(wire_254), .out3(wire_269), .out4(), .out5(), .out6(), .out7());
  TC_Splitter16 # (.UUID(64'd2261501443814513651 ^ UUID)) Splitter16_24 (.in(wire_25[15:0]), .out0(wire_78), .out1());
  TC_Splitter8 # (.UUID(64'd2576232014769382965 ^ UUID)) Splitter8_25 (.in(wire_78), .out0(wire_262), .out1(wire_187), .out2(wire_251), .out3(wire_223), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd2608661849516270155 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_26 (.en(wire_50), .in(wire_132), .out(wire_44_4));
  TC_Switch # (.UUID(64'd746143341221514145 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_27 (.en(wire_18), .in(wire_132), .out(wire_16_2));
  TC_Switch # (.UUID(64'd2038162143482139082 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_28 (.en(wire_75), .in(wire_141), .out(wire_44_2));
  TC_Switch # (.UUID(64'd4451929975376370007 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_29 (.en(wire_8), .in(wire_141), .out(wire_16_0));
  TC_Switch # (.UUID(64'd2149760867058136119 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_30 (.en(wire_106), .in(wire_33), .out(wire_44_0));
  TC_Switch # (.UUID(64'd1120920137235279511 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_31 (.en(wire_88), .in(wire_33), .out(wire_16_1));
  TC_Switch # (.UUID(64'd1049077220225763239 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_32 (.en(wire_36), .in(wire_147), .out(wire_44_1));
  TC_Switch # (.UUID(64'd690331529650965982 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_33 (.en(wire_139), .in(wire_147), .out(wire_16_3));
  TC_Switch # (.UUID(64'd4446234359163774586 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_34 (.en(wire_179), .in(wire_161), .out(wire_44_3));
  TC_Switch # (.UUID(64'd68561501764135042 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_35 (.en(wire_61), .in(wire_161), .out(wire_16_5));
  TC_Switch # (.UUID(64'd2300663947791505692 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_36 (.en(wire_38), .in(wire_86), .out(wire_44_5));
  TC_Switch # (.UUID(64'd1809390294038489791 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_37 (.en(wire_142), .in(wire_86), .out(wire_16_6));
  TC_Switch # (.UUID(64'd2131531128077507626 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_38 (.en(wire_165), .in(wire_138), .out(wire_44_7));
  TC_Switch # (.UUID(64'd2315389642693555300 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_39 (.en(wire_42), .in(wire_138), .out(wire_16_7));
  TC_Switch # (.UUID(64'd4187739606022409523 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_40 (.en(wire_114), .in(wire_214), .out(wire_44_8));
  TC_Switch # (.UUID(64'd1859071114078130426 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_41 (.en(wire_111), .in(wire_214), .out(wire_16_8));
  TC_Equal # (.UUID(64'd137163679941758477 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_42 (.in0(wire_97[15:0]), .in1(wire_156), .out(wire_109));
  TC_Halt # (.UUID(64'd2683931794444888664 ^ UUID)) Halt_43 (.clk(clk), .rst(rst), .en(wire_109));
  TC_Constant # (.UUID(64'd1352990490392554841 ^ UUID), .BIT_WIDTH(64'd16), .value(16'hFFFF)) Constant16_44 (.out(wire_156));
  TC_Switch # (.UUID(64'd971606683869478136 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_45 (.en(wire_103), .in(wire_95[15:0]), .out(wire_44_6));
  TC_Switch # (.UUID(64'd488700789590138722 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_46 (.en(wire_124), .in(wire_13[15:0]), .out(wire_16_4));
  TC_Constant # (.UUID(64'd1219804294531623130 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h0)) Constant16_47 (.out(wire_132));
  TC_Switch # (.UUID(64'd2854432665896608476 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_48 (.en(wire_188), .in(wire_189), .out(wire_260));
  TC_Not # (.UUID(64'd1919204710248089503 ^ UUID), .BIT_WIDTH(64'd1)) Not_49 (.in(wire_109), .out(wire_188));
  TC_Switch # (.UUID(64'd3648642341737646920 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_50 (.en(wire_83), .in(wire_25[15:0]), .out(wire_115));
  TC_Switch # (.UUID(64'd2839537485959427856 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_51 (.en(wire_21), .in(wire_21), .out(wire_83));
  TC_Splitter16 # (.UUID(64'd4451072885120255536 ^ UUID)) Splitter16_52 (.in(wire_97[15:0]), .out0(wire_221), .out1());
  TC_Splitter8 # (.UUID(64'd1191888651688547656 ^ UUID)) Splitter8_53 (.in(wire_221), .out0(wire_129), .out1(wire_37), .out2(wire_224), .out3(wire_219), .out4(), .out5(), .out6(), .out7());
  TC_Not # (.UUID(64'd4189336834672528069 ^ UUID), .BIT_WIDTH(64'd1)) Not_54 (.in(wire_80), .out(wire_118));
  TC_Add # (.UUID(64'd3182557287143411779 ^ UUID), .BIT_WIDTH(64'd16)) Add16_55 (.in0(wire_16), .in1(wire_44), .ci(1'd0), .out(wire_122), .co());
  TC_Add # (.UUID(64'd1424675120960351269 ^ UUID), .BIT_WIDTH(64'd16)) Add16_56 (.in0(wire_16), .in1(wire_25[15:0]), .ci(1'd0), .out(wire_207), .co());
  TC_Switch # (.UUID(64'd284020542177892273 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_57 (.en(wire_119), .in(wire_122), .out(wire_93_0));
  TC_Switch # (.UUID(64'd1034703434088870431 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_58 (.en(wire_53), .in(wire_207), .out(wire_93_1));
  TC_Or # (.UUID(64'd657814780105628035 ^ UUID), .BIT_WIDTH(64'd1)) Or_59 (.in0(wire_21), .in1(wire_53), .out(wire_117));
  TC_Console # (.UUID(64'd1550364046122691923 ^ UUID)) Console_60 (.clk(clk), .rst(rst), .offset({{16{1'b0}}, wire_66 }));
  TC_Ram # (.UUID(64'd2067412014399195219 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd65536)) Ram_61 (.clk(clk), .rst(rst), .load(1'd0), .save(wire_181), .address({{16{1'b0}}, wire_16 }), .in0({{48{1'b0}}, wire_44 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(), .out1(), .out2(), .out3());
  TC_Ram # (.UUID(64'd2804227458846121453 ^ UUID), .WORD_WIDTH(64'd16), .WORD_COUNT(64'd32768)) Ram_62 (.clk(clk), .rst(rst), .load(wire_100), .save(wire_93[0:0]), .address({{16{1'b0}}, wire_44 }), .in0(64'd0), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(), .out1(), .out2(), .out3());
  TC_Splitter16 # (.UUID(64'd763171029710359662 ^ UUID)) Splitter16_63 (.in(wire_93), .out0(), .out1(wire_166));
  TC_Splitter8 # (.UUID(64'd3824024877144842064 ^ UUID)) Splitter8_64 (.in(wire_166), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7(wire_227));
  TC_Decoder1 # (.UUID(64'd4576965811034017994 ^ UUID)) Decoder1_65 (.sel(wire_227), .out0(wire_101), .out1(wire_131));
  TC_Switch # (.UUID(64'd2746301141431459897 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_66 (.en(wire_101), .in(wire_53), .out(wire_235));
  TC_Switch # (.UUID(64'd3430101359472696647 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_67 (.en(wire_101), .in(wire_119), .out(wire_170));
  TC_Switch # (.UUID(64'd1728891745001622010 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_68 (.en(wire_131), .in(wire_119), .out(wire_193));
  TC_Switch # (.UUID(64'd4375680025586519226 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_69 (.en(wire_131), .in(wire_53), .out(wire_100));
  TC_Register # (.UUID(64'd2693553474459199961 ^ UUID), .BIT_WIDTH(64'd16)) Register16_70 (.clk(clk), .rst(rst), .load(wire_77), .save(wire_56), .in(wire_256), .out(wire_66));
  TC_Add # (.UUID(64'd3809269893433252203 ^ UUID), .BIT_WIDTH(64'd16)) Add16_71 (.in0(wire_66), .in1(wire_148), .ci(1'd0), .out(wire_256), .co());
  TC_Constant # (.UUID(64'd2151188605745524424 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_72 (.out(wire_77));
  TC_Constant # (.UUID(64'd1918094738540249611 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h50)) Constant16_73 (.out(wire_148));
  TC_Splitter16 # (.UUID(64'd4494426812884145071 ^ UUID)) Splitter16_74 (.in(wire_97[15:0]), .out0(wire_278), .out1());
  TC_Splitter8 # (.UUID(64'd1684985711211094078 ^ UUID)) Splitter8_75 (.in(wire_278), .out0(wire_281), .out1(wire_94), .out2(wire_247), .out3(wire_19), .out4(), .out5(), .out6(), .out7());
  TC_Not # (.UUID(64'd2891551810552540629 ^ UUID), .BIT_WIDTH(64'd1)) Not_76 (.in(wire_48), .out(wire_250));
  TC_Register # (.UUID(64'd3266843945445956355 ^ UUID), .BIT_WIDTH(64'd16)) Register16_77 (.clk(clk), .rst(rst), .load(wire_266), .save(wire_236), .in(wire_26[15:0]), .out(wire_243));
  TC_Register # (.UUID(64'd373441705232759894 ^ UUID), .BIT_WIDTH(64'd16)) Register16_78 (.clk(clk), .rst(rst), .load(wire_267), .save(wire_123), .in(wire_26[15:0]), .out(wire_158));
  TC_Register # (.UUID(64'd898762616312898673 ^ UUID), .BIT_WIDTH(64'd16)) Register16_79 (.clk(clk), .rst(rst), .load(wire_259), .save(wire_140), .in(wire_26[15:0]), .out(wire_209));
  TC_Register # (.UUID(64'd35259159018310512 ^ UUID), .BIT_WIDTH(64'd16)) Register16_80 (.clk(clk), .rst(rst), .load(wire_121), .save(wire_175), .in(wire_26[15:0]), .out(wire_171));
  TC_Or # (.UUID(64'd3408749404784824565 ^ UUID), .BIT_WIDTH(64'd1)) Or_81 (.in0(wire_63), .in1(wire_159), .out(wire_266));
  TC_Or # (.UUID(64'd2045434085000650231 ^ UUID), .BIT_WIDTH(64'd1)) Or_82 (.in0(wire_2), .in1(wire_152), .out(wire_267));
  TC_Or # (.UUID(64'd4235778316917593708 ^ UUID), .BIT_WIDTH(64'd1)) Or_83 (.in0(wire_199), .in1(wire_160), .out(wire_259));
  TC_Or # (.UUID(64'd1881922342948910945 ^ UUID), .BIT_WIDTH(64'd1)) Or_84 (.in0(wire_39), .in1(wire_49), .out(wire_121));
  TC_Switch # (.UUID(64'd3154836780073834162 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_85 (.en(wire_159), .in(wire_243), .out(wire_44_9));
  TC_Switch # (.UUID(64'd3206739131565530044 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_86 (.en(wire_63), .in(wire_243), .out(wire_16_9));
  TC_Switch # (.UUID(64'd1476550871400967823 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_87 (.en(wire_152), .in(wire_158), .out(wire_44_10));
  TC_Switch # (.UUID(64'd1622071797847061869 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_88 (.en(wire_2), .in(wire_158), .out(wire_16_10));
  TC_Switch # (.UUID(64'd189967047438908968 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_89 (.en(wire_160), .in(wire_209), .out(wire_44_11));
  TC_Switch # (.UUID(64'd3142169352616083849 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_90 (.en(wire_199), .in(wire_209), .out(wire_16_11));
  TC_Switch # (.UUID(64'd2790449206563351533 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_91 (.en(wire_49), .in(wire_171), .out(wire_44_12));
  TC_Switch # (.UUID(64'd1382504743536358321 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_92 (.en(wire_39), .in(wire_171), .out(wire_16_12));
  TC_DotMatrixDisplay # (.UUID(64'd2660535027850879501 ^ UUID)) DotMatrixDisplay_93 (.clk(clk), .rst(rst), .en_y(wire_24[0:0]), .en_x(wire_20[0:0]), .color_info(wire_24[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd1287415170352733091 ^ UUID)) DotMatrixDisplay_94 (.clk(clk), .rst(rst), .en_y(wire_9[0:0]), .en_x(wire_20[0:0]), .color_info(wire_9[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd4375632836552484410 ^ UUID)) DotMatrixDisplay_95 (.clk(clk), .rst(rst), .en_y(wire_51[0:0]), .en_x(wire_20[0:0]), .color_info(wire_51[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd4352128498737539568 ^ UUID)) DotMatrixDisplay_96 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_20[0:0]), .color_info(wire_17[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd4375805759909017124 ^ UUID)) DotMatrixDisplay_97 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_20[0:0]), .color_info(wire_22[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd4001708814053949966 ^ UUID)) DotMatrixDisplay_98 (.clk(clk), .rst(rst), .en_y(wire_31[0:0]), .en_x(wire_20[0:0]), .color_info(wire_31[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd3789421783879759989 ^ UUID)) DotMatrixDisplay_99 (.clk(clk), .rst(rst), .en_y(wire_59[0:0]), .en_x(wire_20[0:0]), .color_info(wire_59[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd3949917514357280402 ^ UUID)) DotMatrixDisplay_100 (.clk(clk), .rst(rst), .en_y(wire_58[0:0]), .en_x(wire_64[0:0]), .color_info(wire_58[31:0]), .pixel_info(wire_64));
  TC_DotMatrixDisplay # (.UUID(64'd1120366264718111392 ^ UUID)) DotMatrixDisplay_101 (.clk(clk), .rst(rst), .en_y(wire_24[0:0]), .en_x(wire_64[0:0]), .color_info(wire_24[31:0]), .pixel_info(wire_64));
  TC_DotMatrixDisplay # (.UUID(64'd3830190475406040627 ^ UUID)) DotMatrixDisplay_102 (.clk(clk), .rst(rst), .en_y(wire_9[0:0]), .en_x(wire_64[0:0]), .color_info(wire_9[31:0]), .pixel_info(wire_64));
  TC_DotMatrixDisplay # (.UUID(64'd3695649649918959220 ^ UUID)) DotMatrixDisplay_103 (.clk(clk), .rst(rst), .en_y(wire_51[0:0]), .en_x(wire_64[0:0]), .color_info(wire_51[31:0]), .pixel_info(wire_64));
  TC_DotMatrixDisplay # (.UUID(64'd2190167902128485018 ^ UUID)) DotMatrixDisplay_104 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_64[0:0]), .color_info(wire_17[31:0]), .pixel_info(wire_64));
  TC_DotMatrixDisplay # (.UUID(64'd108023444932811778 ^ UUID)) DotMatrixDisplay_105 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_10[0:0]), .color_info(wire_17[31:0]), .pixel_info(wire_10));
  TC_DotMatrixDisplay # (.UUID(64'd3127548314519555293 ^ UUID)) DotMatrixDisplay_106 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_64[0:0]), .color_info(wire_22[31:0]), .pixel_info(wire_64));
  TC_DotMatrixDisplay # (.UUID(64'd3232957164641830670 ^ UUID)) DotMatrixDisplay_107 (.clk(clk), .rst(rst), .en_y(wire_59[0:0]), .en_x(wire_64[0:0]), .color_info(wire_59[31:0]), .pixel_info(wire_64));
  TC_DotMatrixDisplay # (.UUID(64'd2013870924499775536 ^ UUID)) DotMatrixDisplay_108 (.clk(clk), .rst(rst), .en_y(wire_58[0:0]), .en_x(wire_10[0:0]), .color_info(wire_58[31:0]), .pixel_info(wire_10));
  TC_DotMatrixDisplay # (.UUID(64'd1700230642759998846 ^ UUID)) DotMatrixDisplay_109 (.clk(clk), .rst(rst), .en_y(wire_24[0:0]), .en_x(wire_10[0:0]), .color_info(wire_24[31:0]), .pixel_info(wire_10));
  TC_DotMatrixDisplay # (.UUID(64'd640862205653523348 ^ UUID)) DotMatrixDisplay_110 (.clk(clk), .rst(rst), .en_y(wire_9[0:0]), .en_x(wire_10[0:0]), .color_info(wire_9[31:0]), .pixel_info(wire_10));
  TC_DotMatrixDisplay # (.UUID(64'd1441056504049384023 ^ UUID)) DotMatrixDisplay_111 (.clk(clk), .rst(rst), .en_y(wire_51[0:0]), .en_x(wire_10[0:0]), .color_info(wire_51[31:0]), .pixel_info(wire_10));
  TC_DotMatrixDisplay # (.UUID(64'd4360991051994526462 ^ UUID)) DotMatrixDisplay_112 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_40[0:0]), .color_info(wire_17[31:0]), .pixel_info(wire_40));
  TC_DotMatrixDisplay # (.UUID(64'd3732720467344721449 ^ UUID)) DotMatrixDisplay_113 (.clk(clk), .rst(rst), .en_y(wire_31[0:0]), .en_x(wire_64[0:0]), .color_info(wire_31[31:0]), .pixel_info(wire_64));
  TC_DotMatrixDisplay # (.UUID(64'd3164120181411694497 ^ UUID)) DotMatrixDisplay_114 (.clk(clk), .rst(rst), .en_y(wire_31[0:0]), .en_x(wire_10[0:0]), .color_info(wire_31[31:0]), .pixel_info(wire_10));
  TC_DotMatrixDisplay # (.UUID(64'd3058994005473620099 ^ UUID)) DotMatrixDisplay_115 (.clk(clk), .rst(rst), .en_y(wire_59[0:0]), .en_x(wire_10[0:0]), .color_info(wire_59[31:0]), .pixel_info(wire_10));
  TC_DotMatrixDisplay # (.UUID(64'd3043865689462340485 ^ UUID)) DotMatrixDisplay_116 (.clk(clk), .rst(rst), .en_y(wire_58[0:0]), .en_x(wire_40[0:0]), .color_info(wire_58[31:0]), .pixel_info(wire_40));
  TC_DotMatrixDisplay # (.UUID(64'd1232256408208860842 ^ UUID)) DotMatrixDisplay_117 (.clk(clk), .rst(rst), .en_y(wire_24[0:0]), .en_x(wire_40[0:0]), .color_info(wire_24[31:0]), .pixel_info(wire_40));
  TC_DotMatrixDisplay # (.UUID(64'd456775015865694566 ^ UUID)) DotMatrixDisplay_118 (.clk(clk), .rst(rst), .en_y(wire_9[0:0]), .en_x(wire_40[0:0]), .color_info(wire_9[31:0]), .pixel_info(wire_40));
  TC_DotMatrixDisplay # (.UUID(64'd1486947349792475943 ^ UUID)) DotMatrixDisplay_119 (.clk(clk), .rst(rst), .en_y(wire_51[0:0]), .en_x(wire_40[0:0]), .color_info(wire_51[31:0]), .pixel_info(wire_40));
  TC_DotMatrixDisplay # (.UUID(64'd1986390658814520529 ^ UUID)) DotMatrixDisplay_120 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_10[0:0]), .color_info(wire_22[31:0]), .pixel_info(wire_10));
  TC_DotMatrixDisplay # (.UUID(64'd428599916565265934 ^ UUID)) DotMatrixDisplay_121 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_40[0:0]), .color_info(wire_22[31:0]), .pixel_info(wire_40));
  TC_DotMatrixDisplay # (.UUID(64'd1361741769374930265 ^ UUID)) DotMatrixDisplay_122 (.clk(clk), .rst(rst), .en_y(wire_31[0:0]), .en_x(wire_40[0:0]), .color_info(wire_31[31:0]), .pixel_info(wire_40));
  TC_DotMatrixDisplay # (.UUID(64'd3810902491231665649 ^ UUID)) DotMatrixDisplay_123 (.clk(clk), .rst(rst), .en_y(wire_59[0:0]), .en_x(wire_40[0:0]), .color_info(wire_59[31:0]), .pixel_info(wire_40));
  TC_DotMatrixDisplay # (.UUID(64'd145789043302394905 ^ UUID)) DotMatrixDisplay_124 (.clk(clk), .rst(rst), .en_y(wire_58[0:0]), .en_x(wire_43[0:0]), .color_info(wire_58[31:0]), .pixel_info(wire_43));
  TC_DotMatrixDisplay # (.UUID(64'd3780736919653097053 ^ UUID)) DotMatrixDisplay_125 (.clk(clk), .rst(rst), .en_y(wire_24[0:0]), .en_x(wire_43[0:0]), .color_info(wire_24[31:0]), .pixel_info(wire_43));
  TC_DotMatrixDisplay # (.UUID(64'd2485800408185936591 ^ UUID)) DotMatrixDisplay_126 (.clk(clk), .rst(rst), .en_y(wire_9[0:0]), .en_x(wire_43[0:0]), .color_info(wire_9[31:0]), .pixel_info(wire_43));
  TC_DotMatrixDisplay # (.UUID(64'd3637982062020866444 ^ UUID)) DotMatrixDisplay_127 (.clk(clk), .rst(rst), .en_y(wire_51[0:0]), .en_x(wire_43[0:0]), .color_info(wire_51[31:0]), .pixel_info(wire_43));
  TC_DotMatrixDisplay # (.UUID(64'd2077992963286351604 ^ UUID)) DotMatrixDisplay_128 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_43[0:0]), .color_info(wire_17[31:0]), .pixel_info(wire_43));
  TC_DotMatrixDisplay # (.UUID(64'd3780255053339576859 ^ UUID)) DotMatrixDisplay_129 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_43[0:0]), .color_info(wire_22[31:0]), .pixel_info(wire_43));
  TC_DotMatrixDisplay # (.UUID(64'd3088612785393467744 ^ UUID)) DotMatrixDisplay_130 (.clk(clk), .rst(rst), .en_y(wire_31[0:0]), .en_x(wire_43[0:0]), .color_info(wire_31[31:0]), .pixel_info(wire_43));
  TC_DotMatrixDisplay # (.UUID(64'd4340287621202113208 ^ UUID)) DotMatrixDisplay_131 (.clk(clk), .rst(rst), .en_y(wire_59[0:0]), .en_x(wire_43[0:0]), .color_info(wire_59[31:0]), .pixel_info(wire_43));
  TC_DotMatrixDisplay # (.UUID(64'd3263142337545802511 ^ UUID)) DotMatrixDisplay_132 (.clk(clk), .rst(rst), .en_y(wire_58[0:0]), .en_x(wire_0[0:0]), .color_info(wire_58[31:0]), .pixel_info(wire_0));
  TC_DotMatrixDisplay # (.UUID(64'd4368304585025255821 ^ UUID)) DotMatrixDisplay_133 (.clk(clk), .rst(rst), .en_y(wire_24[0:0]), .en_x(wire_0[0:0]), .color_info(wire_24[31:0]), .pixel_info(wire_0));
  TC_DotMatrixDisplay # (.UUID(64'd3035154864325599620 ^ UUID)) DotMatrixDisplay_134 (.clk(clk), .rst(rst), .en_y(wire_9[0:0]), .en_x(wire_0[0:0]), .color_info(wire_9[31:0]), .pixel_info(wire_0));
  TC_DotMatrixDisplay # (.UUID(64'd1984067145119237049 ^ UUID)) DotMatrixDisplay_135 (.clk(clk), .rst(rst), .en_y(wire_51[0:0]), .en_x(wire_0[0:0]), .color_info(wire_51[31:0]), .pixel_info(wire_0));
  TC_DotMatrixDisplay # (.UUID(64'd257903097512365689 ^ UUID)) DotMatrixDisplay_136 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_0[0:0]), .color_info(wire_17[31:0]), .pixel_info(wire_0));
  TC_DotMatrixDisplay # (.UUID(64'd1855803350615582069 ^ UUID)) DotMatrixDisplay_137 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_0[0:0]), .color_info(wire_22[31:0]), .pixel_info(wire_0));
  TC_DotMatrixDisplay # (.UUID(64'd4156190447566119276 ^ UUID)) DotMatrixDisplay_138 (.clk(clk), .rst(rst), .en_y(wire_31[0:0]), .en_x(wire_0[0:0]), .color_info(wire_31[31:0]), .pixel_info(wire_0));
  TC_DotMatrixDisplay # (.UUID(64'd3549196530068966916 ^ UUID)) DotMatrixDisplay_139 (.clk(clk), .rst(rst), .en_y(wire_59[0:0]), .en_x(wire_0[0:0]), .color_info(wire_59[31:0]), .pixel_info(wire_0));
  TC_DotMatrixDisplay # (.UUID(64'd3746276803240527606 ^ UUID)) DotMatrixDisplay_140 (.clk(clk), .rst(rst), .en_y(wire_58[0:0]), .en_x(wire_20[0:0]), .color_info(wire_58[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd4237472817339994162 ^ UUID)) DotMatrixDisplay_141 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_20[0:0]), .color_info(wire_92[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd1177830180225486220 ^ UUID)) DotMatrixDisplay_142 (.clk(clk), .rst(rst), .en_y(wire_12[0:0]), .en_x(wire_20[0:0]), .color_info(wire_12[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd250680188831281298 ^ UUID)) DotMatrixDisplay_143 (.clk(clk), .rst(rst), .en_y(wire_5[0:0]), .en_x(wire_20[0:0]), .color_info(wire_5[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd1576462328986410349 ^ UUID)) DotMatrixDisplay_144 (.clk(clk), .rst(rst), .en_y(wire_27[0:0]), .en_x(wire_20[0:0]), .color_info(wire_27[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd316625153349409673 ^ UUID)) DotMatrixDisplay_145 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_20[0:0]), .color_info(wire_102[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd959143668139620378 ^ UUID)) DotMatrixDisplay_146 (.clk(clk), .rst(rst), .en_y(wire_28[0:0]), .en_x(wire_20[0:0]), .color_info(wire_28[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd684938010714015909 ^ UUID)) DotMatrixDisplay_147 (.clk(clk), .rst(rst), .en_y(wire_52[0:0]), .en_x(wire_20[0:0]), .color_info(wire_52[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd1796769576252909689 ^ UUID)) DotMatrixDisplay_148 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_64[0:0]), .color_info(wire_23[31:0]), .pixel_info(wire_64));
  TC_DotMatrixDisplay # (.UUID(64'd28266181691657389 ^ UUID)) DotMatrixDisplay_149 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_64[0:0]), .color_info(wire_92[31:0]), .pixel_info(wire_64));
  TC_DotMatrixDisplay # (.UUID(64'd3196962412568546329 ^ UUID)) DotMatrixDisplay_150 (.clk(clk), .rst(rst), .en_y(wire_12[0:0]), .en_x(wire_64[0:0]), .color_info(wire_12[31:0]), .pixel_info(wire_64));
  TC_DotMatrixDisplay # (.UUID(64'd2205871638966640606 ^ UUID)) DotMatrixDisplay_151 (.clk(clk), .rst(rst), .en_y(wire_5[0:0]), .en_x(wire_64[0:0]), .color_info(wire_5[31:0]), .pixel_info(wire_64));
  TC_DotMatrixDisplay # (.UUID(64'd3874186372446959361 ^ UUID)) DotMatrixDisplay_152 (.clk(clk), .rst(rst), .en_y(wire_27[0:0]), .en_x(wire_64[0:0]), .color_info(wire_27[31:0]), .pixel_info(wire_64));
  TC_DotMatrixDisplay # (.UUID(64'd2720360903878823189 ^ UUID)) DotMatrixDisplay_153 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_64[0:0]), .color_info(wire_102[31:0]), .pixel_info(wire_64));
  TC_DotMatrixDisplay # (.UUID(64'd504346027738870704 ^ UUID)) DotMatrixDisplay_154 (.clk(clk), .rst(rst), .en_y(wire_28[0:0]), .en_x(wire_64[0:0]), .color_info(wire_28[31:0]), .pixel_info(wire_64));
  TC_DotMatrixDisplay # (.UUID(64'd184655924988308158 ^ UUID)) DotMatrixDisplay_155 (.clk(clk), .rst(rst), .en_y(wire_52[0:0]), .en_x(wire_64[0:0]), .color_info(wire_52[31:0]), .pixel_info(wire_64));
  TC_DotMatrixDisplay # (.UUID(64'd3162126675592577790 ^ UUID)) DotMatrixDisplay_156 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_10[0:0]), .color_info(wire_23[31:0]), .pixel_info(wire_10));
  TC_DotMatrixDisplay # (.UUID(64'd841957664227372441 ^ UUID)) DotMatrixDisplay_157 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_10[0:0]), .color_info(wire_92[31:0]), .pixel_info(wire_10));
  TC_DotMatrixDisplay # (.UUID(64'd4388146087367304388 ^ UUID)) DotMatrixDisplay_158 (.clk(clk), .rst(rst), .en_y(wire_12[0:0]), .en_x(wire_10[0:0]), .color_info(wire_12[31:0]), .pixel_info(wire_10));
  TC_DotMatrixDisplay # (.UUID(64'd935756330229132165 ^ UUID)) DotMatrixDisplay_159 (.clk(clk), .rst(rst), .en_y(wire_5[0:0]), .en_x(wire_10[0:0]), .color_info(wire_5[31:0]), .pixel_info(wire_10));
  TC_DotMatrixDisplay # (.UUID(64'd38018604794773973 ^ UUID)) DotMatrixDisplay_160 (.clk(clk), .rst(rst), .en_y(wire_27[0:0]), .en_x(wire_10[0:0]), .color_info(wire_27[31:0]), .pixel_info(wire_10));
  TC_DotMatrixDisplay # (.UUID(64'd1334297701942639290 ^ UUID)) DotMatrixDisplay_161 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_10[0:0]), .color_info(wire_102[31:0]), .pixel_info(wire_10));
  TC_DotMatrixDisplay # (.UUID(64'd971239419644370685 ^ UUID)) DotMatrixDisplay_162 (.clk(clk), .rst(rst), .en_y(wire_28[0:0]), .en_x(wire_10[0:0]), .color_info(wire_28[31:0]), .pixel_info(wire_10));
  TC_DotMatrixDisplay # (.UUID(64'd2299276613863097833 ^ UUID)) DotMatrixDisplay_163 (.clk(clk), .rst(rst), .en_y(wire_52[0:0]), .en_x(wire_10[0:0]), .color_info(wire_52[31:0]), .pixel_info(wire_10));
  TC_DotMatrixDisplay # (.UUID(64'd4066308585007913895 ^ UUID)) DotMatrixDisplay_164 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_40[0:0]), .color_info(wire_23[31:0]), .pixel_info(wire_40));
  TC_DotMatrixDisplay # (.UUID(64'd1188730429928185190 ^ UUID)) DotMatrixDisplay_165 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_40[0:0]), .color_info(wire_92[31:0]), .pixel_info(wire_40));
  TC_DotMatrixDisplay # (.UUID(64'd4280800355417676313 ^ UUID)) DotMatrixDisplay_166 (.clk(clk), .rst(rst), .en_y(wire_12[0:0]), .en_x(wire_40[0:0]), .color_info(wire_12[31:0]), .pixel_info(wire_40));
  TC_DotMatrixDisplay # (.UUID(64'd4360520332522264149 ^ UUID)) DotMatrixDisplay_167 (.clk(clk), .rst(rst), .en_y(wire_5[0:0]), .en_x(wire_40[0:0]), .color_info(wire_5[31:0]), .pixel_info(wire_40));
  TC_DotMatrixDisplay # (.UUID(64'd475575386071264203 ^ UUID)) DotMatrixDisplay_168 (.clk(clk), .rst(rst), .en_y(wire_27[0:0]), .en_x(wire_40[0:0]), .color_info(wire_27[31:0]), .pixel_info(wire_40));
  TC_DotMatrixDisplay # (.UUID(64'd4099921249160036118 ^ UUID)) DotMatrixDisplay_169 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_40[0:0]), .color_info(wire_102[31:0]), .pixel_info(wire_40));
  TC_DotMatrixDisplay # (.UUID(64'd2008157871612466016 ^ UUID)) DotMatrixDisplay_170 (.clk(clk), .rst(rst), .en_y(wire_28[0:0]), .en_x(wire_40[0:0]), .color_info(wire_28[31:0]), .pixel_info(wire_40));
  TC_DotMatrixDisplay # (.UUID(64'd3526081255155773975 ^ UUID)) DotMatrixDisplay_171 (.clk(clk), .rst(rst), .en_y(wire_52[0:0]), .en_x(wire_40[0:0]), .color_info(wire_52[31:0]), .pixel_info(wire_40));
  TC_DotMatrixDisplay # (.UUID(64'd1085763782026657154 ^ UUID)) DotMatrixDisplay_172 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_43[0:0]), .color_info(wire_23[31:0]), .pixel_info(wire_43));
  TC_DotMatrixDisplay # (.UUID(64'd1935004646604641077 ^ UUID)) DotMatrixDisplay_173 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_43[0:0]), .color_info(wire_92[31:0]), .pixel_info(wire_43));
  TC_DotMatrixDisplay # (.UUID(64'd4228153944513970773 ^ UUID)) DotMatrixDisplay_174 (.clk(clk), .rst(rst), .en_y(wire_12[0:0]), .en_x(wire_43[0:0]), .color_info(wire_12[31:0]), .pixel_info(wire_43));
  TC_DotMatrixDisplay # (.UUID(64'd3380853135653261586 ^ UUID)) DotMatrixDisplay_175 (.clk(clk), .rst(rst), .en_y(wire_5[0:0]), .en_x(wire_43[0:0]), .color_info(wire_5[31:0]), .pixel_info(wire_43));
  TC_DotMatrixDisplay # (.UUID(64'd142464094186867413 ^ UUID)) DotMatrixDisplay_176 (.clk(clk), .rst(rst), .en_y(wire_27[0:0]), .en_x(wire_43[0:0]), .color_info(wire_27[31:0]), .pixel_info(wire_43));
  TC_DotMatrixDisplay # (.UUID(64'd988217888803392985 ^ UUID)) DotMatrixDisplay_177 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_43[0:0]), .color_info(wire_102[31:0]), .pixel_info(wire_43));
  TC_DotMatrixDisplay # (.UUID(64'd54720530278277779 ^ UUID)) DotMatrixDisplay_178 (.clk(clk), .rst(rst), .en_y(wire_28[0:0]), .en_x(wire_43[0:0]), .color_info(wire_28[31:0]), .pixel_info(wire_43));
  TC_DotMatrixDisplay # (.UUID(64'd2688678971804628028 ^ UUID)) DotMatrixDisplay_179 (.clk(clk), .rst(rst), .en_y(wire_52[0:0]), .en_x(wire_43[0:0]), .color_info(wire_52[31:0]), .pixel_info(wire_43));
  TC_DotMatrixDisplay # (.UUID(64'd553058778145918310 ^ UUID)) DotMatrixDisplay_180 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_0[0:0]), .color_info(wire_23[31:0]), .pixel_info(wire_0));
  TC_DotMatrixDisplay # (.UUID(64'd2098597773896322169 ^ UUID)) DotMatrixDisplay_181 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_0[0:0]), .color_info(wire_92[31:0]), .pixel_info(wire_0));
  TC_DotMatrixDisplay # (.UUID(64'd1919740307961683958 ^ UUID)) DotMatrixDisplay_182 (.clk(clk), .rst(rst), .en_y(wire_12[0:0]), .en_x(wire_0[0:0]), .color_info(wire_12[31:0]), .pixel_info(wire_0));
  TC_DotMatrixDisplay # (.UUID(64'd2955390637246533656 ^ UUID)) DotMatrixDisplay_183 (.clk(clk), .rst(rst), .en_y(wire_5[0:0]), .en_x(wire_0[0:0]), .color_info(wire_5[31:0]), .pixel_info(wire_0));
  TC_DotMatrixDisplay # (.UUID(64'd3399628396733223633 ^ UUID)) DotMatrixDisplay_184 (.clk(clk), .rst(rst), .en_y(wire_27[0:0]), .en_x(wire_0[0:0]), .color_info(wire_27[31:0]), .pixel_info(wire_0));
  TC_DotMatrixDisplay # (.UUID(64'd1503255611657110166 ^ UUID)) DotMatrixDisplay_185 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_0[0:0]), .color_info(wire_102[31:0]), .pixel_info(wire_0));
  TC_DotMatrixDisplay # (.UUID(64'd1934210770642016723 ^ UUID)) DotMatrixDisplay_186 (.clk(clk), .rst(rst), .en_y(wire_28[0:0]), .en_x(wire_0[0:0]), .color_info(wire_28[31:0]), .pixel_info(wire_0));
  TC_DotMatrixDisplay # (.UUID(64'd4430890296674284431 ^ UUID)) DotMatrixDisplay_187 (.clk(clk), .rst(rst), .en_y(wire_52[0:0]), .en_x(wire_0[0:0]), .color_info(wire_52[31:0]), .pixel_info(wire_0));
  TC_DotMatrixDisplay # (.UUID(64'd1370192036403734636 ^ UUID)) DotMatrixDisplay_188 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_20[0:0]), .color_info(wire_23[31:0]), .pixel_info(wire_20));
  TC_DotMatrixDisplay # (.UUID(64'd1914293527285665104 ^ UUID)) DotMatrixDisplay_189 (.clk(clk), .rst(rst), .en_y(wire_58[0:0]), .en_x(wire_14[0:0]), .color_info(wire_58[31:0]), .pixel_info(wire_14));
  TC_DotMatrixDisplay # (.UUID(64'd4024378624965788820 ^ UUID)) DotMatrixDisplay_190 (.clk(clk), .rst(rst), .en_y(wire_24[0:0]), .en_x(wire_14[0:0]), .color_info(wire_24[31:0]), .pixel_info(wire_14));
  TC_DotMatrixDisplay # (.UUID(64'd331796838499445221 ^ UUID)) DotMatrixDisplay_191 (.clk(clk), .rst(rst), .en_y(wire_9[0:0]), .en_x(wire_14[0:0]), .color_info(wire_9[31:0]), .pixel_info(wire_14));
  TC_DotMatrixDisplay # (.UUID(64'd1109146203016946320 ^ UUID)) DotMatrixDisplay_192 (.clk(clk), .rst(rst), .en_y(wire_51[0:0]), .en_x(wire_14[0:0]), .color_info(wire_51[31:0]), .pixel_info(wire_14));
  TC_DotMatrixDisplay # (.UUID(64'd2037862037394616530 ^ UUID)) DotMatrixDisplay_193 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_14[0:0]), .color_info(wire_17[31:0]), .pixel_info(wire_14));
  TC_DotMatrixDisplay # (.UUID(64'd756317346051932726 ^ UUID)) DotMatrixDisplay_194 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_14[0:0]), .color_info(wire_22[31:0]), .pixel_info(wire_14));
  TC_DotMatrixDisplay # (.UUID(64'd741221856880638315 ^ UUID)) DotMatrixDisplay_195 (.clk(clk), .rst(rst), .en_y(wire_31[0:0]), .en_x(wire_14[0:0]), .color_info(wire_31[31:0]), .pixel_info(wire_14));
  TC_DotMatrixDisplay # (.UUID(64'd2554897745454830451 ^ UUID)) DotMatrixDisplay_196 (.clk(clk), .rst(rst), .en_y(wire_59[0:0]), .en_x(wire_14[0:0]), .color_info(wire_59[31:0]), .pixel_info(wire_14));
  TC_DotMatrixDisplay # (.UUID(64'd4352234980297914729 ^ UUID)) DotMatrixDisplay_197 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_14[0:0]), .color_info(wire_23[31:0]), .pixel_info(wire_14));
  TC_DotMatrixDisplay # (.UUID(64'd4044674900922762564 ^ UUID)) DotMatrixDisplay_198 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_14[0:0]), .color_info(wire_92[31:0]), .pixel_info(wire_14));
  TC_DotMatrixDisplay # (.UUID(64'd2175572511635428388 ^ UUID)) DotMatrixDisplay_199 (.clk(clk), .rst(rst), .en_y(wire_12[0:0]), .en_x(wire_14[0:0]), .color_info(wire_12[31:0]), .pixel_info(wire_14));
  TC_DotMatrixDisplay # (.UUID(64'd1352766524066348872 ^ UUID)) DotMatrixDisplay_200 (.clk(clk), .rst(rst), .en_y(wire_5[0:0]), .en_x(wire_14[0:0]), .color_info(wire_5[31:0]), .pixel_info(wire_14));
  TC_DotMatrixDisplay # (.UUID(64'd1625039672493008527 ^ UUID)) DotMatrixDisplay_201 (.clk(clk), .rst(rst), .en_y(wire_27[0:0]), .en_x(wire_14[0:0]), .color_info(wire_27[31:0]), .pixel_info(wire_14));
  TC_DotMatrixDisplay # (.UUID(64'd672361543425103183 ^ UUID)) DotMatrixDisplay_202 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_14[0:0]), .color_info(wire_102[31:0]), .pixel_info(wire_14));
  TC_DotMatrixDisplay # (.UUID(64'd1607234245481583786 ^ UUID)) DotMatrixDisplay_203 (.clk(clk), .rst(rst), .en_y(wire_28[0:0]), .en_x(wire_14[0:0]), .color_info(wire_28[31:0]), .pixel_info(wire_14));
  TC_DotMatrixDisplay # (.UUID(64'd2377050978244241774 ^ UUID)) DotMatrixDisplay_204 (.clk(clk), .rst(rst), .en_y(wire_52[0:0]), .en_x(wire_14[0:0]), .color_info(wire_52[31:0]), .pixel_info(wire_14));
  TC_DotMatrixDisplay # (.UUID(64'd3222873545553085433 ^ UUID)) DotMatrixDisplay_205 (.clk(clk), .rst(rst), .en_y(wire_58[0:0]), .en_x(wire_68[0:0]), .color_info(wire_58[31:0]), .pixel_info(wire_68));
  TC_DotMatrixDisplay # (.UUID(64'd3188765738163086443 ^ UUID)) DotMatrixDisplay_206 (.clk(clk), .rst(rst), .en_y(wire_24[0:0]), .en_x(wire_68[0:0]), .color_info(wire_24[31:0]), .pixel_info(wire_68));
  TC_DotMatrixDisplay # (.UUID(64'd838700140978907233 ^ UUID)) DotMatrixDisplay_207 (.clk(clk), .rst(rst), .en_y(wire_9[0:0]), .en_x(wire_68[0:0]), .color_info(wire_9[31:0]), .pixel_info(wire_68));
  TC_DotMatrixDisplay # (.UUID(64'd3920730297055212015 ^ UUID)) DotMatrixDisplay_208 (.clk(clk), .rst(rst), .en_y(wire_51[0:0]), .en_x(wire_68[0:0]), .color_info(wire_51[31:0]), .pixel_info(wire_68));
  TC_DotMatrixDisplay # (.UUID(64'd3481948759443637 ^ UUID)) DotMatrixDisplay_209 (.clk(clk), .rst(rst), .en_y(wire_17[0:0]), .en_x(wire_68[0:0]), .color_info(wire_17[31:0]), .pixel_info(wire_68));
  TC_DotMatrixDisplay # (.UUID(64'd511172518486640794 ^ UUID)) DotMatrixDisplay_210 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_68[0:0]), .color_info(wire_22[31:0]), .pixel_info(wire_68));
  TC_DotMatrixDisplay # (.UUID(64'd4053020964562097569 ^ UUID)) DotMatrixDisplay_211 (.clk(clk), .rst(rst), .en_y(wire_31[0:0]), .en_x(wire_68[0:0]), .color_info(wire_31[31:0]), .pixel_info(wire_68));
  TC_DotMatrixDisplay # (.UUID(64'd3303805443456392646 ^ UUID)) DotMatrixDisplay_212 (.clk(clk), .rst(rst), .en_y(wire_59[0:0]), .en_x(wire_68[0:0]), .color_info(wire_59[31:0]), .pixel_info(wire_68));
  TC_DotMatrixDisplay # (.UUID(64'd3229541704842781328 ^ UUID)) DotMatrixDisplay_213 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_68[0:0]), .color_info(wire_23[31:0]), .pixel_info(wire_68));
  TC_DotMatrixDisplay # (.UUID(64'd1520258463232062736 ^ UUID)) DotMatrixDisplay_214 (.clk(clk), .rst(rst), .en_y(wire_92[0:0]), .en_x(wire_68[0:0]), .color_info(wire_92[31:0]), .pixel_info(wire_68));
  TC_DotMatrixDisplay # (.UUID(64'd3535073739167951615 ^ UUID)) DotMatrixDisplay_215 (.clk(clk), .rst(rst), .en_y(wire_12[0:0]), .en_x(wire_68[0:0]), .color_info(wire_12[31:0]), .pixel_info(wire_68));
  TC_DotMatrixDisplay # (.UUID(64'd2508590195121546232 ^ UUID)) DotMatrixDisplay_216 (.clk(clk), .rst(rst), .en_y(wire_5[0:0]), .en_x(wire_68[0:0]), .color_info(wire_5[31:0]), .pixel_info(wire_68));
  TC_DotMatrixDisplay # (.UUID(64'd4190156087276806644 ^ UUID)) DotMatrixDisplay_217 (.clk(clk), .rst(rst), .en_y(wire_27[0:0]), .en_x(wire_68[0:0]), .color_info(wire_27[31:0]), .pixel_info(wire_68));
  TC_DotMatrixDisplay # (.UUID(64'd3357160141127693591 ^ UUID)) DotMatrixDisplay_218 (.clk(clk), .rst(rst), .en_y(wire_102[0:0]), .en_x(wire_68[0:0]), .color_info(wire_102[31:0]), .pixel_info(wire_68));
  TC_DotMatrixDisplay # (.UUID(64'd3712829154125709738 ^ UUID)) DotMatrixDisplay_219 (.clk(clk), .rst(rst), .en_y(wire_28[0:0]), .en_x(wire_68[0:0]), .color_info(wire_28[31:0]), .pixel_info(wire_68));
  TC_DotMatrixDisplay # (.UUID(64'd2545725033216246256 ^ UUID)) DotMatrixDisplay_220 (.clk(clk), .rst(rst), .en_y(wire_52[0:0]), .en_x(wire_68[0:0]), .color_info(wire_52[31:0]), .pixel_info(wire_68));
  TC_Mul # (.UUID(64'd2748524405844472327 ^ UUID), .BIT_WIDTH(64'd16)) DivMod16_221 (.in0(wire_44), .in1(wire_81), .out0(wire_35), .out1(wire_99));
  TC_Mul # (.UUID(64'd4020347048163863131 ^ UUID), .BIT_WIDTH(64'd16)) DivMod16_222 (.in0(wire_16), .in1(wire_195), .out0(wire_212), .out1(wire_127));
  TC_Constant # (.UUID(64'd1313141643564538265 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h6)) Constant16_223 (.out(wire_195));
  TC_Constant # (.UUID(64'd4112089032370153264 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h8)) Constant16_224 (.out(wire_81));
  TC_Splitter16 # (.UUID(64'd2668786745693159507 ^ UUID)) Splitter16_225 (.in(wire_212), .out0(wire_135), .out1());
  TC_Splitter8 # (.UUID(64'd2631886754935636255 ^ UUID)) Splitter8_226 (.in(wire_135), .out0(wire_226), .out1(wire_264), .out2(wire_220), .out3(wire_268), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd550414518326034956 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_227 (.en(wire_7), .in(wire_32), .out(wire_58));
  TC_Switch # (.UUID(64'd977382900955430648 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_228 (.en(wire_162), .in(wire_32), .out(wire_24));
  TC_Switch # (.UUID(64'd1891242292111482311 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_229 (.en(wire_167), .in(wire_32), .out(wire_9));
  TC_Switch # (.UUID(64'd856889246029500943 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_230 (.en(wire_110), .in(wire_32), .out(wire_51));
  TC_Switch # (.UUID(64'd3189954206832060770 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_231 (.en(wire_1), .in(wire_32), .out(wire_17));
  TC_Switch # (.UUID(64'd2600416908798528202 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_232 (.en(wire_144), .in(wire_32), .out(wire_22));
  TC_Switch # (.UUID(64'd3352059561228947819 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_233 (.en(wire_85), .in(wire_32), .out(wire_31));
  TC_Switch # (.UUID(64'd3576546926653500711 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_234 (.en(wire_237), .in(wire_32), .out(wire_59));
  TC_Switch # (.UUID(64'd773945265408688934 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_235 (.en(wire_105), .in(wire_32), .out(wire_23));
  TC_Switch # (.UUID(64'd4124677947420211807 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_236 (.en(wire_151), .in(wire_32), .out(wire_92));
  TC_Switch # (.UUID(64'd1892597805610563739 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_237 (.en(wire_164), .in(wire_32), .out(wire_12));
  TC_Switch # (.UUID(64'd4501036839557111240 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_238 (.en(wire_180), .in(wire_32), .out(wire_5));
  TC_Switch # (.UUID(64'd2653282250793028984 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_239 (.en(wire_55), .in(wire_32), .out(wire_27));
  TC_Switch # (.UUID(64'd2835551167096927095 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_240 (.en(wire_82), .in(wire_32), .out(wire_102));
  TC_Switch # (.UUID(64'd811538821685340963 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_241 (.en(wire_67), .in(wire_32), .out(wire_28));
  TC_Switch # (.UUID(64'd1795419328706358879 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_242 (.en(wire_41), .in(wire_32), .out(wire_52));
  TC_Switch # (.UUID(64'd3384031002647223712 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_243 (.en(wire_65), .in(wire_62), .out(wire_20));
  TC_Switch # (.UUID(64'd796360369331162321 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_244 (.en(wire_248), .in(wire_62), .out(wire_64));
  TC_Switch # (.UUID(64'd770893388854325356 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_245 (.en(wire_125), .in(wire_62), .out(wire_10));
  TC_Switch # (.UUID(64'd2296729005521048932 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_246 (.en(wire_104), .in(wire_62), .out(wire_40));
  TC_Switch # (.UUID(64'd2700874401252926434 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_247 (.en(wire_11), .in(wire_62), .out(wire_43));
  TC_Switch # (.UUID(64'd3871697537247032043 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_248 (.en(wire_242), .in(wire_62), .out(wire_0));
  TC_Switch # (.UUID(64'd1657382633537052929 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_249 (.en(wire_194), .in(wire_62), .out(wire_14));
  TC_Switch # (.UUID(64'd2430440528996199989 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_250 (.en(wire_87), .in(wire_62), .out(wire_68));
  TC_Splitter8 # (.UUID(64'd4038412651713004570 ^ UUID)) Splitter8_251 (.in(wire_261), .out0(wire_47), .out1(wire_96), .out2(wire_137), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter16 # (.UUID(64'd3776431078096079195 ^ UUID)) Splitter16_252 (.in(wire_35), .out0(wire_261), .out1());
  TC_Decoder3 # (.UUID(64'd4013734321313478962 ^ UUID)) Decoder3_253 (.dis(wire_204), .sel0(wire_47), .sel1(wire_96), .sel2(wire_137), .out0(wire_182), .out1(wire_178), .out2(wire_275), .out3(wire_172), .out4(wire_203), .out5(wire_3), .out6(wire_69), .out7(wire_246));
  TC_Maker64 # (.UUID(64'd1192448886920089561 ^ UUID)) Maker64_254 (.in0(wire_155), .in1(wire_253), .in2(wire_232), .in3(wire_206), .in4(8'd0), .in5(8'd0), .in6(8'd0), .in7(8'd0), .out(wire_32));
  TC_Mux # (.UUID(64'd3182122184138242733 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_255 (.sel(wire_29), .in0(wire_222), .in1(wire_184), .out(wire_62));
  TC_Constant # (.UUID(64'd499839709284412840 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_256 (.out(wire_155));
  TC_Register # (.UUID(64'd3760785338326490848 ^ UUID), .BIT_WIDTH(64'd8)) Register8_257 (.clk(clk), .rst(rst), .load(wire_6), .save(wire_57), .in(wire_79), .out(wire_206));
  TC_Register # (.UUID(64'd4329544050407358966 ^ UUID), .BIT_WIDTH(64'd8)) Register8_258 (.clk(clk), .rst(rst), .load(wire_6), .save(wire_57), .in(wire_169), .out(wire_232));
  TC_Register # (.UUID(64'd199054775600590363 ^ UUID), .BIT_WIDTH(64'd8)) Register8_259 (.clk(clk), .rst(rst), .load(wire_6), .save(wire_57), .in(wire_168), .out(wire_253));
  TC_Constant # (.UUID(64'd224588895404758285 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_260 (.out(wire_6));
  TC_Splitter16 # (.UUID(64'd2025205086175333323 ^ UUID)) Splitter16_261 (.in(wire_16), .out0(wire_79), .out1(wire_169));
  TC_Splitter16 # (.UUID(64'd2367030245059056516 ^ UUID)) Splitter16_262 (.in(wire_44), .out0(wire_168), .out1());
  TC_Constant # (.UUID(64'd1704767967961521854 ^ UUID), .BIT_WIDTH(64'd64), .value(64'h0)) Constant64_263 (.out(wire_222));
  TC_Not # (.UUID(64'd1573479007334595178 ^ UUID), .BIT_WIDTH(64'd1)) Not_264 (.in(wire_89), .out(wire_215));
  TC_Not # (.UUID(64'd4448026403053823646 ^ UUID), .BIT_WIDTH(64'd1)) Not_265 (.in(wire_89), .out(wire_204));
  TC_Maker64 # (.UUID(64'd509307949451829158 ^ UUID)) Maker64_266 (.in0(wire_280), .in1(wire_190), .in2(wire_91), .in3(wire_197), .in4(wire_258), .in5(wire_183), .in6(wire_113), .in7(wire_225), .out(wire_192));
  TC_Switch # (.UUID(64'd3450977581660059279 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_267 (.en(wire_112), .in(wire_84), .out(wire_190));
  TC_Switch # (.UUID(64'd3243380833679066833 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_268 (.en(wire_202), .in(wire_84), .out(wire_91));
  TC_Switch # (.UUID(64'd1815840084729226412 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_269 (.en(wire_228), .in(wire_84), .out(wire_197));
  TC_Switch # (.UUID(64'd4246131709043477595 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_270 (.en(wire_149), .in(wire_84), .out(wire_258));
  TC_Switch # (.UUID(64'd3003808122831947155 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_271 (.en(wire_30), .in(wire_84), .out(wire_183));
  TC_Switch # (.UUID(64'd573612594436248865 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_272 (.en(wire_108), .in(wire_84), .out(wire_113));
  TC_Constant # (.UUID(64'd3268609550269517760 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_273 (.out(wire_280));
  TC_Constant # (.UUID(64'd1513805053441976731 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_274 (.out(wire_225));
  TC_Maker8 # (.UUID(64'd2761932721413399018 ^ UUID)) Maker8_275 (.in0(wire_255), .in1(wire_208), .in2(wire_201), .in3(wire_116), .in4(wire_213), .in5(wire_90), .in6(wire_218), .in7(wire_177), .out(wire_84));
  TC_Decoder3 # (.UUID(64'd2669229198398327855 ^ UUID)) Decoder3_276 (.dis(wire_71), .sel0(wire_233), .sel1(wire_249), .sel2(wire_274), .out0(wire_112), .out1(wire_202), .out2(wire_228), .out3(wire_149), .out4(wire_30), .out5(wire_108), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd2415290327339560914 ^ UUID)) Decoder3_277 (.dis(wire_71), .sel0(wire_154), .sel1(wire_272), .sel2(wire_238), .out0(wire_174), .out1(wire_210), .out2(wire_273), .out3(wire_263), .out4(wire_234), .out5(wire_196), .out6(wire_231), .out7(wire_60));
  TC_Splitter8 # (.UUID(64'd4390030900946952921 ^ UUID)) Splitter8_278 (.in(wire_127[7:0]), .out0(wire_233), .out1(wire_249), .out2(wire_274), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd3413845568106834524 ^ UUID)) Splitter8_279 (.in(wire_99[7:0]), .out0(wire_154), .out1(wire_272), .out2(wire_238), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Not # (.UUID(64'd2354531697599582148 ^ UUID), .BIT_WIDTH(64'd1)) Not_280 (.in(wire_89), .out(wire_71));
  OPP8 # (.UUID(64'd1987821792969644964 ^ UUID)) OPP8_281 (.clk(clk), .rst(rst), .Input_1(wire_182), .Input_2(wire_178), .Input_3(wire_275), .Input_4(wire_172), .Input_5(wire_203), .Input_6(wire_3), .Input_7(wire_69), .Input_8(wire_246), .Enable_All(wire_72), .Output_1(wire_65), .Output_2(wire_248), .Output_3(wire_125), .Output_4(wire_104), .Output_5(wire_11), .Output_6(wire_242), .Output_7(wire_194), .Output_8(wire_87));
  OPP16 # (.UUID(64'd2240121763827152286 ^ UUID)) OPP16_282 (.clk(clk), .rst(rst), .Input_1(wire_257), .Input_2(wire_217), .Input_3(wire_186), .Input_4(wire_229), .Input_5(wire_241), .Input_6(wire_211), .Input_7(wire_153), .Input_8(wire_270), .Input_9(wire_198), .Input_10(wire_252), .Input_11(wire_271), .Input_12(wire_143), .Input_13(wire_4), .Input_14(wire_107), .Input_15(wire_46), .Input_16(wire_200), .Enable_All(wire_72), .Output_1(wire_41), .Output_2(wire_67), .Output_3(wire_82), .Output_4(wire_55), .Output_5(wire_180), .Output_6(wire_164), .Output_7(wire_151), .Output_8(wire_105), .Output_9(wire_237), .Output_10(wire_85), .Output_11(wire_144), .Output_12(wire_1), .Output_13(wire_110), .Output_14(wire_167), .Output_15(wire_162), .Output_16(wire_7));
  OPP8 # (.UUID(64'd511775211755439032 ^ UUID)) OPP8_283 (.clk(clk), .rst(rst), .Input_1(wire_174), .Input_2(wire_210), .Input_3(wire_273), .Input_4(wire_263), .Input_5(wire_234), .Input_6(wire_196), .Input_7(wire_231), .Input_8(wire_60), .Enable_All(1'd0), .Output_1(wire_255), .Output_2(wire_208), .Output_3(wire_201), .Output_4(wire_116), .Output_5(wire_213), .Output_6(wire_90), .Output_7(wire_218), .Output_8(wire_177));
  DEC2 # (.UUID(64'd771286428991844547 ^ UUID)) DEC2_284 (.clk(clk), .rst(rst), .Input_1(wire_240), .Input_2(wire_176), .Disable(wire_109), .Output_1(wire_45), .Output_2(wire_80), .Output_3(wire_48), .Output_4(wire_15));
  DEC4 # (.UUID(64'd971863642718444548 ^ UUID)) DEC4_285 (.clk(clk), .rst(rst), .Bit_1(wire_130), .Bit_2(wire_185), .Bit_3(wire_239), .Bit_4(wire_277), .Disable(wire_124), .Output_1(wire_142), .Output_2(wire_42), .Output_3(wire_111), .Output_4(wire_61), .Output_5(wire_139), .Output_6(wire_88), .Output_7(wire_8), .Output_8(wire_18), .Output_9(wire_63), .Output_10(wire_2), .Output_11(wire_199), .Output_12(wire_39), .Output_13(), .Output_14(), .Output_15(), .Output_16());
  DEC4 # (.UUID(64'd1590120432676397143 ^ UUID)) DEC4_286 (.clk(clk), .rst(rst), .Bit_1(wire_216), .Bit_2(wire_98), .Bit_3(wire_254), .Bit_4(wire_269), .Disable(wire_103), .Output_1(wire_38), .Output_2(wire_165), .Output_3(wire_114), .Output_4(wire_179), .Output_5(wire_36), .Output_6(wire_106), .Output_7(wire_75), .Output_8(wire_50), .Output_9(wire_159), .Output_10(wire_152), .Output_11(wire_160), .Output_12(wire_49), .Output_13(), .Output_14(), .Output_15(), .Output_16());
  DEC4 # (.UUID(64'd3642349192148398088 ^ UUID)) DEC4_287 (.clk(clk), .rst(rst), .Bit_1(wire_262), .Bit_2(wire_187), .Bit_3(wire_251), .Bit_4(wire_223), .Disable(wire_117), .Output_1(wire_73), .Output_2(wire_34), .Output_3(wire_74), .Output_4(wire_136), .Output_5(wire_70), .Output_6(wire_205), .Output_7(wire_150), .Output_8(wire_145), .Output_9(wire_236), .Output_10(wire_123), .Output_11(wire_140), .Output_12(wire_175), .Output_13(), .Output_14(), .Output_15(), .Output_16());
  DEC4 # (.UUID(64'd4338106330534265481 ^ UUID)) DEC4_288 (.clk(clk), .rst(rst), .Bit_1(wire_281), .Bit_2(wire_94), .Bit_3(wire_247), .Bit_4(wire_19), .Disable(wire_250), .Output_1(wire_146), .Output_2(wire_54), .Output_3(), .Output_4(wire_72), .Output_5(wire_57), .Output_6(wire_89), .Output_7(wire_56), .Output_8(wire_181), .Output_9(), .Output_10(), .Output_11(), .Output_12(), .Output_13(), .Output_14(), .Output_15(), .Output_16());
  DEC4 # (.UUID(64'd2116072289912876009 ^ UUID)) DEC4_289 (.clk(clk), .rst(rst), .Bit_1(wire_129), .Bit_2(wire_37), .Bit_3(wire_224), .Bit_4(wire_219), .Disable(wire_118), .Output_1(), .Output_2(), .Output_3(), .Output_4(), .Output_5(), .Output_6(), .Output_7(wire_53), .Output_8(wire_119), .Output_9(), .Output_10(), .Output_11(), .Output_12(), .Output_13(), .Output_14(), .Output_15(), .Output_16());
  DEC4 # (.UUID(64'd2389694038429158952 ^ UUID)) DEC4_290 (.clk(clk), .rst(rst), .Bit_1(wire_226), .Bit_2(wire_264), .Bit_3(wire_220), .Bit_4(wire_268), .Disable(wire_215), .Output_1(wire_211), .Output_2(wire_153), .Output_3(wire_270), .Output_4(wire_241), .Output_5(wire_229), .Output_6(wire_186), .Output_7(wire_217), .Output_8(wire_257), .Output_9(wire_198), .Output_10(wire_252), .Output_11(wire_271), .Output_12(wire_143), .Output_13(wire_4), .Output_14(wire_107), .Output_15(wire_46), .Output_16(wire_200));
  ALU # (.UUID(64'd2633888247542289904 ^ UUID)) ALU_291 (.clk(clk), .rst(rst), .Instruction(wire_97[15:0]), .Input_1(wire_16), .Input_2(wire_44), .Enable(wire_15), .Output(wire_26_1[15:0]));
  COND # (.UUID(64'd1460830942441319647 ^ UUID)) COND_292 (.clk(clk), .rst(rst), .Instruction(wire_97[15:0]), .Input_1(wire_16), .Input_2(wire_44), .Enable(wire_45), .Output(wire_21));
  TC_Mux # (.UUID(64'd1000091076309775908 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_293 (.sel(wire_72), .in0(wire_192), .in1(wire_76), .out(wire_184));
  TC_Constant # (.UUID(64'd2073010886631854991 ^ UUID), .BIT_WIDTH(64'd64), .value(64'h1FFFFFFFFFFFF01)) Constant64_294 (.out(wire_76));
  TC_Or # (.UUID(64'd2275862259491790157 ^ UUID), .BIT_WIDTH(64'd1)) Or_295 (.in0(wire_89), .in1(wire_72), .out(wire_29));
  TC_Switch # (.UUID(64'd4021291688878439030 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_296 (.en(wire_54), .in(wire_244), .out(wire_26_3[7:0]));
  TC_Switch # (.UUID(64'd4156448496845195677 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_297 (.en(wire_133), .in({{7{1'b0}}, wire_134 }), .out(wire_244));
  TC_Switch # (.UUID(64'd3594967734502713487 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_298 (.en(wire_146), .in({{7{1'b0}}, wire_276 }), .out(wire_26_2[7:0]));

  wire [63:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [63:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [63:0] wire_9;
  wire [63:0] wire_10;
  wire [0:0] wire_11;
  wire [63:0] wire_12;
  wire [63:0] wire_13;
  wire [63:0] wire_14;
  wire [0:0] wire_15;
  wire [15:0] wire_16;
  wire [15:0] wire_16_0;
  wire [15:0] wire_16_1;
  wire [15:0] wire_16_2;
  wire [15:0] wire_16_3;
  wire [15:0] wire_16_4;
  wire [15:0] wire_16_5;
  wire [15:0] wire_16_6;
  wire [15:0] wire_16_7;
  wire [15:0] wire_16_8;
  wire [15:0] wire_16_9;
  wire [15:0] wire_16_10;
  wire [15:0] wire_16_11;
  wire [15:0] wire_16_12;
  assign wire_16 = wire_16_0|wire_16_1|wire_16_2|wire_16_3|wire_16_4|wire_16_5|wire_16_6|wire_16_7|wire_16_8|wire_16_9|wire_16_10|wire_16_11|wire_16_12;
  wire [63:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [63:0] wire_20;
  wire [0:0] wire_21;
  wire [63:0] wire_22;
  wire [63:0] wire_23;
  wire [63:0] wire_24;
  wire [63:0] wire_25;
  wire [63:0] wire_26;
  wire [63:0] wire_26_0;
  wire [63:0] wire_26_1;
  wire [63:0] wire_26_2;
  wire [63:0] wire_26_3;
  assign wire_26 = wire_26_0|wire_26_1|wire_26_2|wire_26_3;
  wire [63:0] wire_27;
  wire [63:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [63:0] wire_31;
  wire [63:0] wire_32;
  wire [15:0] wire_33;
  wire [0:0] wire_34;
  wire [15:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [63:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [63:0] wire_43;
  wire [15:0] wire_44;
  wire [15:0] wire_44_0;
  wire [15:0] wire_44_1;
  wire [15:0] wire_44_2;
  wire [15:0] wire_44_3;
  wire [15:0] wire_44_4;
  wire [15:0] wire_44_5;
  wire [15:0] wire_44_6;
  wire [15:0] wire_44_7;
  wire [15:0] wire_44_8;
  wire [15:0] wire_44_9;
  wire [15:0] wire_44_10;
  wire [15:0] wire_44_11;
  wire [15:0] wire_44_12;
  assign wire_44 = wire_44_0|wire_44_1|wire_44_2|wire_44_3|wire_44_4|wire_44_5|wire_44_6|wire_44_7|wire_44_8|wire_44_9|wire_44_10|wire_44_11|wire_44_12;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [63:0] wire_51;
  wire [63:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [63:0] wire_58;
  wire [63:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [63:0] wire_62;
  wire [0:0] wire_63;
  wire [63:0] wire_64;
  wire [0:0] wire_65;
  wire [15:0] wire_66;
  wire [0:0] wire_67;
  wire [63:0] wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [0:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [63:0] wire_76;
  wire [0:0] wire_77;
  wire [7:0] wire_78;
  wire [7:0] wire_79;
  wire [0:0] wire_80;
  wire [15:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;
  wire [7:0] wire_84;
  wire [0:0] wire_85;
  wire [15:0] wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;
  wire [0:0] wire_90;
  wire [7:0] wire_91;
  wire [63:0] wire_92;
  wire [15:0] wire_93;
  wire [15:0] wire_93_0;
  wire [15:0] wire_93_1;
  assign wire_93 = wire_93_0|wire_93_1;
  wire [0:0] wire_94;
  wire [63:0] wire_95;
  wire [0:0] wire_96;
  wire [63:0] wire_97;
  wire [0:0] wire_98;
  wire [15:0] wire_99;
  wire [0:0] wire_100;
  wire [0:0] wire_101;
  wire [63:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [0:0] wire_105;
  wire [0:0] wire_106;
  wire [0:0] wire_107;
  wire [0:0] wire_108;
  wire [0:0] wire_109;
  wire [0:0] wire_110;
  wire [0:0] wire_111;
  wire [0:0] wire_112;
  wire [7:0] wire_113;
  wire [0:0] wire_114;
  wire [15:0] wire_115;
  wire [0:0] wire_116;
  wire [0:0] wire_117;
  wire [0:0] wire_118;
  wire [0:0] wire_119;
  wire [0:0] wire_120;
  wire [0:0] wire_121;
  wire [15:0] wire_122;
  wire [0:0] wire_123;
  wire [0:0] wire_124;
  wire [0:0] wire_125;
  wire [15:0] wire_126;
  wire [15:0] wire_127;
  wire [0:0] wire_128;
  wire [0:0] wire_129;
  wire [0:0] wire_130;
  wire [0:0] wire_131;
  wire [15:0] wire_132;
  wire [0:0] wire_133;
  assign wire_133 = 0;
  wire [0:0] wire_134;
  assign wire_134 = 0;
  wire [7:0] wire_135;
  wire [0:0] wire_136;
  wire [0:0] wire_137;
  wire [15:0] wire_138;
  wire [0:0] wire_139;
  wire [0:0] wire_140;
  wire [15:0] wire_141;
  wire [0:0] wire_142;
  wire [0:0] wire_143;
  wire [0:0] wire_144;
  wire [0:0] wire_145;
  wire [0:0] wire_146;
  wire [15:0] wire_147;
  wire [15:0] wire_148;
  wire [0:0] wire_149;
  wire [0:0] wire_150;
  wire [0:0] wire_151;
  wire [0:0] wire_152;
  wire [0:0] wire_153;
  wire [0:0] wire_154;
  wire [7:0] wire_155;
  wire [15:0] wire_156;
  wire [7:0] wire_157;
  wire [15:0] wire_158;
  wire [0:0] wire_159;
  wire [0:0] wire_160;
  wire [15:0] wire_161;
  wire [0:0] wire_162;
  wire [0:0] wire_163;
  wire [0:0] wire_164;
  wire [0:0] wire_165;
  wire [7:0] wire_166;
  wire [0:0] wire_167;
  wire [7:0] wire_168;
  wire [7:0] wire_169;
  wire [0:0] wire_170;
  wire [15:0] wire_171;
  wire [0:0] wire_172;
  wire [0:0] wire_173;
  wire [0:0] wire_174;
  wire [0:0] wire_175;
  wire [0:0] wire_176;
  wire [0:0] wire_177;
  wire [0:0] wire_178;
  wire [0:0] wire_179;
  wire [0:0] wire_180;
  wire [0:0] wire_181;
  wire [0:0] wire_182;
  wire [7:0] wire_183;
  wire [63:0] wire_184;
  wire [0:0] wire_185;
  wire [0:0] wire_186;
  wire [0:0] wire_187;
  wire [0:0] wire_188;
  wire [7:0] wire_189;
  wire [7:0] wire_190;
  wire [7:0] wire_191;
  wire [63:0] wire_192;
  wire [0:0] wire_193;
  wire [0:0] wire_194;
  wire [15:0] wire_195;
  wire [0:0] wire_196;
  wire [7:0] wire_197;
  wire [0:0] wire_198;
  wire [0:0] wire_199;
  wire [0:0] wire_200;
  wire [0:0] wire_201;
  wire [0:0] wire_202;
  wire [0:0] wire_203;
  wire [0:0] wire_204;
  wire [0:0] wire_205;
  wire [7:0] wire_206;
  wire [15:0] wire_207;
  wire [0:0] wire_208;
  wire [15:0] wire_209;
  wire [0:0] wire_210;
  wire [0:0] wire_211;
  wire [15:0] wire_212;
  wire [0:0] wire_213;
  wire [15:0] wire_214;
  wire [0:0] wire_215;
  wire [0:0] wire_216;
  wire [0:0] wire_217;
  wire [0:0] wire_218;
  wire [0:0] wire_219;
  wire [0:0] wire_220;
  wire [7:0] wire_221;
  wire [63:0] wire_222;
  wire [0:0] wire_223;
  wire [0:0] wire_224;
  wire [7:0] wire_225;
  wire [0:0] wire_226;
  wire [0:0] wire_227;
  wire [0:0] wire_228;
  wire [0:0] wire_229;
  wire [0:0] wire_230;
  wire [0:0] wire_231;
  wire [7:0] wire_232;
  wire [0:0] wire_233;
  wire [0:0] wire_234;
  wire [0:0] wire_235;
  wire [0:0] wire_236;
  wire [0:0] wire_237;
  wire [0:0] wire_238;
  wire [0:0] wire_239;
  wire [0:0] wire_240;
  wire [0:0] wire_241;
  wire [0:0] wire_242;
  wire [15:0] wire_243;
  wire [7:0] wire_244;
  wire [0:0] wire_245;
  wire [0:0] wire_246;
  wire [0:0] wire_247;
  wire [0:0] wire_248;
  wire [0:0] wire_249;
  wire [0:0] wire_250;
  wire [0:0] wire_251;
  wire [0:0] wire_252;
  wire [7:0] wire_253;
  wire [0:0] wire_254;
  wire [0:0] wire_255;
  wire [15:0] wire_256;
  wire [0:0] wire_257;
  wire [7:0] wire_258;
  wire [0:0] wire_259;
  wire [7:0] wire_260;
  wire [7:0] wire_261;
  wire [0:0] wire_262;
  wire [0:0] wire_263;
  wire [0:0] wire_264;
  wire [0:0] wire_265;
  wire [0:0] wire_266;
  wire [0:0] wire_267;
  wire [0:0] wire_268;
  wire [0:0] wire_269;
  wire [0:0] wire_270;
  wire [0:0] wire_271;
  wire [0:0] wire_272;
  wire [0:0] wire_273;
  wire [0:0] wire_274;
  wire [0:0] wire_275;
  wire [0:0] wire_276;
  assign wire_276 = 0;
  wire [0:0] wire_277;
  wire [7:0] wire_278;
  wire [0:0] wire_279;
  wire [7:0] wire_280;
  wire [0:0] wire_281;

endmodule
