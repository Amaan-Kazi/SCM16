module DEC4 (clk, rst, Bit_1, Bit_2, Bit_3, Bit_4, Disable, Output_1, Output_2, Output_3, Output_4, Output_5, Output_6, Output_7, Output_8, Output_9, Output_10, Output_11, Output_12, Output_13, Output_14, Output_15, Output_16);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] Bit_1;
  input  wire [0:0] Bit_2;
  input  wire [0:0] Bit_3;
  input  wire [0:0] Bit_4;
  input  wire [0:0] Disable;
  output  wire [0:0] Output_1;
  output  wire [0:0] Output_2;
  output  wire [0:0] Output_3;
  output  wire [0:0] Output_4;
  output  wire [0:0] Output_5;
  output  wire [0:0] Output_6;
  output  wire [0:0] Output_7;
  output  wire [0:0] Output_8;
  output  wire [0:0] Output_9;
  output  wire [0:0] Output_10;
  output  wire [0:0] Output_11;
  output  wire [0:0] Output_12;
  output  wire [0:0] Output_13;
  output  wire [0:0] Output_14;
  output  wire [0:0] Output_15;
  output  wire [0:0] Output_16;

  TC_Decoder3 # (.UUID(64'd2265727218055464636 ^ UUID)) Decoder3_0 (.dis(wire_22), .sel0(wire_8), .sel1(wire_7), .sel2(wire_15), .out0(wire_23), .out1(wire_12), .out2(wire_16), .out3(wire_11), .out4(wire_21), .out5(wire_9), .out6(wire_5), .out7(wire_2));
  TC_Decoder3 # (.UUID(64'd4151446233815205602 ^ UUID)) Decoder3_1 (.dis(wire_10), .sel0(wire_8), .sel1(wire_7), .sel2(wire_15), .out0(wire_17), .out1(wire_13), .out2(wire_1), .out3(wire_14), .out4(wire_19), .out5(wire_6), .out6(wire_20), .out7(wire_3));
  TC_Or # (.UUID(64'd1144441976216115803 ^ UUID), .BIT_WIDTH(64'd1)) Or_2 (.in0(wire_4), .in1(wire_0), .out(wire_22));
  TC_Or # (.UUID(64'd1448808864368720956 ^ UUID), .BIT_WIDTH(64'd1)) Or_3 (.in0(wire_4), .in1(wire_18), .out(wire_10));
  TC_Not # (.UUID(64'd1948449524954060999 ^ UUID), .BIT_WIDTH(64'd1)) Not_4 (.in(wire_0), .out(wire_18));
  TC_Splitter8 # (.UUID(64'd2392041343466285091 ^ UUID)) Splitter8_5 (.in(8'd0), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd2955497353746114555 ^ UUID)) Splitter8_6 (.in(8'd0), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd1586858191449826786 ^ UUID)) Splitter8_7 (.in(8'd0), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd1420095608691041084 ^ UUID)) Splitter8_8 (.in(8'd0), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd484362997219790821 ^ UUID)) Splitter8_9 (.in(8'd0), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd2845739053448873615 ^ UUID)) Splitter8_10 (.in(8'd0), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd937364978927028657 ^ UUID)) Splitter8_11 (.in(8'd0), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd3238714810038928330 ^ UUID)) Splitter8_12 (.in(8'd0), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7());

  wire [0:0] wire_0;
  assign wire_0 = Bit_4;
  wire [0:0] wire_1;
  assign Output_11 = wire_1;
  wire [0:0] wire_2;
  assign Output_3 = wire_2;
  wire [0:0] wire_3;
  assign Output_16 = wire_3;
  wire [0:0] wire_4;
  assign wire_4 = Disable;
  wire [0:0] wire_5;
  assign Output_2 = wire_5;
  wire [0:0] wire_6;
  assign Output_14 = wire_6;
  wire [0:0] wire_7;
  assign wire_7 = Bit_2;
  wire [0:0] wire_8;
  assign wire_8 = Bit_1;
  wire [0:0] wire_9;
  assign Output_1 = wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  assign Output_5 = wire_11;
  wire [0:0] wire_12;
  assign Output_7 = wire_12;
  wire [0:0] wire_13;
  assign Output_10 = wire_13;
  wire [0:0] wire_14;
  assign Output_12 = wire_14;
  wire [0:0] wire_15;
  assign wire_15 = Bit_3;
  wire [0:0] wire_16;
  assign Output_6 = wire_16;
  wire [0:0] wire_17;
  assign Output_9 = wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  assign Output_13 = wire_19;
  wire [0:0] wire_20;
  assign Output_15 = wire_20;
  wire [0:0] wire_21;
  assign Output_4 = wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  assign Output_8 = wire_23;

endmodule
