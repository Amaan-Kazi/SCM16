module SCM16 (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_Program # (.UUID(64'd3036675205634735936 ^ UUID), .WORD_WIDTH(64'd16), .DEFAULT_FILE_NAME("Program_2A247002B2183F40.w16.bin"), .ARG_SIG("Program_2A247002B2183F40=%s")) Program_0 (.clk(clk), .rst(rst), .address(wire_126), .out0(wire_18), .out1(wire_59), .out2(wire_19), .out3(wire_2));
  TC_Counter # (.UUID(64'd3613463651816973605 ^ UUID), .BIT_WIDTH(64'd16), .count(16'd4)) Counter16_1 (.clk(clk), .rst(rst), .save(wire_8), .in(wire_63), .out(wire_126));
  TC_Ram # (.UUID(64'd3779316721177258366 ^ UUID), .WORD_WIDTH(64'd16), .WORD_COUNT(64'd32768)) Ram_2 (.clk(clk), .rst(rst), .load(wire_81), .save(wire_113), .address({{16{1'b0}}, wire_1 }), .in0({{48{1'b0}}, wire_15 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_30_1), .out1(), .out2(), .out3());
  TC_Splitter16 # (.UUID(64'd1964885700083813915 ^ UUID)) Splitter16_3 (.in(wire_18[15:0]), .out0(), .out1(wire_127));
  TC_Splitter8 # (.UUID(64'd2865909427779811686 ^ UUID)) Splitter8_4 (.in(wire_121), .out0(), .out1(), .out2(), .out3(), .out4(wire_125), .out5(wire_44), .out6(wire_46), .out7(wire_73));
  TC_Register # (.UUID(64'd1768297580719965166 ^ UUID), .BIT_WIDTH(64'd16)) Register16_5 (.clk(clk), .rst(rst), .load(wire_35), .save(wire_56), .in(wire_30[15:0]), .out(wire_21));
  TC_Register # (.UUID(64'd12270441446668041 ^ UUID), .BIT_WIDTH(64'd16)) Register16_6 (.clk(clk), .rst(rst), .load(wire_92), .save(wire_41), .in(wire_30[15:0]), .out(wire_98));
  TC_Register # (.UUID(64'd3602252881066521773 ^ UUID), .BIT_WIDTH(64'd16)) Register16_7 (.clk(clk), .rst(rst), .load(wire_105), .save(wire_16), .in(wire_30[15:0]), .out(wire_17));
  TC_Register # (.UUID(64'd937036284257795972 ^ UUID), .BIT_WIDTH(64'd16)) Register16_8 (.clk(clk), .rst(rst), .load(wire_110), .save(wire_20), .in(wire_30[15:0]), .out(wire_86));
  TC_Register # (.UUID(64'd1771485704314964723 ^ UUID), .BIT_WIDTH(64'd16)) Register16_9 (.clk(clk), .rst(rst), .load(wire_27), .save(wire_58), .in(wire_30[15:0]), .out(wire_68));
  TC_Register # (.UUID(64'd1030977193978425972 ^ UUID), .BIT_WIDTH(64'd16)) Register16_10 (.clk(clk), .rst(rst), .load(wire_99), .save(wire_42), .in(wire_30[15:0]), .out(wire_76));
  TC_Register # (.UUID(64'd1897207591897939717 ^ UUID), .BIT_WIDTH(64'd16)) Register16_11 (.clk(clk), .rst(rst), .load(wire_50), .save(wire_38), .in(wire_30[15:0]), .out(wire_117));
  TC_Splitter16 # (.UUID(64'd1676756795661497062 ^ UUID)) Splitter16_12 (.in(wire_59[15:0]), .out0(wire_109), .out1());
  TC_Splitter16 # (.UUID(64'd2723123645093883319 ^ UUID)) Splitter16_13 (.in(wire_19[15:0]), .out0(wire_13), .out1());
  TC_Or # (.UUID(64'd3489109707031568152 ^ UUID), .BIT_WIDTH(64'd1)) Or_14 (.in0(wire_64), .in1(wire_43), .out(wire_107));
  TC_Or # (.UUID(64'd2757568662684548394 ^ UUID), .BIT_WIDTH(64'd1)) Or_15 (.in0(wire_97), .in1(wire_80), .out(wire_35));
  TC_Or # (.UUID(64'd2444150779797091056 ^ UUID), .BIT_WIDTH(64'd1)) Or_16 (.in0(wire_88), .in1(wire_11), .out(wire_92));
  TC_Or # (.UUID(64'd3998494940572441480 ^ UUID), .BIT_WIDTH(64'd1)) Or_17 (.in0(wire_55), .in1(wire_9), .out(wire_105));
  TC_Or # (.UUID(64'd3745487864523206918 ^ UUID), .BIT_WIDTH(64'd1)) Or_18 (.in0(wire_23), .in1(wire_22), .out(wire_110));
  TC_Or # (.UUID(64'd151306593792916243 ^ UUID), .BIT_WIDTH(64'd1)) Or_19 (.in0(wire_5), .in1(wire_53), .out(wire_27));
  TC_Or # (.UUID(64'd3493104666195700629 ^ UUID), .BIT_WIDTH(64'd1)) Or_20 (.in0(wire_47), .in1(wire_69), .out(wire_99));
  TC_Or # (.UUID(64'd3870924515638343503 ^ UUID), .BIT_WIDTH(64'd1)) Or_21 (.in0(wire_4), .in1(wire_51), .out(wire_50));
  TC_Splitter8 # (.UUID(64'd2466557324773763251 ^ UUID)) Splitter8_22 (.in(wire_109), .out0(wire_111), .out1(wire_118), .out2(wire_67), .out3(wire_128), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd1977466255751035882 ^ UUID)) Splitter8_23 (.in(wire_13), .out0(wire_60), .out1(wire_114), .out2(wire_79), .out3(wire_71), .out4(), .out5(), .out6(), .out7());
  TC_Splitter16 # (.UUID(64'd2261501443814513651 ^ UUID)) Splitter16_24 (.in(wire_2[15:0]), .out0(wire_87), .out1());
  TC_Splitter8 # (.UUID(64'd2576232014769382965 ^ UUID)) Splitter8_25 (.in(wire_87), .out0(wire_93), .out1(wire_119), .out2(wire_104), .out3(wire_112), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd2608661849516270155 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_26 (.en(wire_43), .in(wire_14), .out(wire_15_11));
  TC_Switch # (.UUID(64'd746143341221514145 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_27 (.en(wire_64), .in(wire_14), .out(wire_24_11));
  TC_Switch # (.UUID(64'd2038162143482139082 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_28 (.en(wire_80), .in(wire_21), .out(wire_15_10));
  TC_Switch # (.UUID(64'd4451929975376370007 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_29 (.en(wire_97), .in(wire_21), .out(wire_24_10));
  TC_Switch # (.UUID(64'd2149760867058136119 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_30 (.en(wire_11), .in(wire_98), .out(wire_15_9));
  TC_Switch # (.UUID(64'd1120920137235279511 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_31 (.en(wire_88), .in(wire_98), .out(wire_24_9));
  TC_Switch # (.UUID(64'd1049077220225763239 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_32 (.en(wire_9), .in(wire_17), .out(wire_15_8));
  TC_Switch # (.UUID(64'd690331529650965982 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_33 (.en(wire_55), .in(wire_17), .out(wire_24_8));
  TC_Switch # (.UUID(64'd4446234359163774586 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_34 (.en(wire_22), .in(wire_86), .out(wire_15_7));
  TC_Switch # (.UUID(64'd68561501764135042 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_35 (.en(wire_23), .in(wire_86), .out(wire_24_7));
  TC_Switch # (.UUID(64'd2300663947791505692 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_36 (.en(wire_53), .in(wire_68), .out(wire_15_5));
  TC_Switch # (.UUID(64'd1809390294038489791 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_37 (.en(wire_5), .in(wire_68), .out(wire_24_6));
  TC_Switch # (.UUID(64'd2131531128077507626 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_38 (.en(wire_69), .in(wire_76), .out(wire_15_3));
  TC_Switch # (.UUID(64'd2315389642693555300 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_39 (.en(wire_47), .in(wire_76), .out(wire_24_5));
  TC_Switch # (.UUID(64'd4187739606022409523 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_40 (.en(wire_51), .in(wire_117), .out(wire_15_1));
  TC_Switch # (.UUID(64'd1859071114078130426 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_41 (.en(wire_4), .in(wire_117), .out(wire_24_4));
  TC_Equal # (.UUID(64'd137163679941758477 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_42 (.in0(wire_18[15:0]), .in1(wire_94), .out(wire_12));
  TC_Halt # (.UUID(64'd2683931794444888664 ^ UUID)) Halt_43 (.clk(clk), .rst(rst), .en(wire_12));
  TC_Constant # (.UUID(64'd1352990490392554841 ^ UUID), .BIT_WIDTH(64'd16), .value(16'hFFFF)) Constant16_44 (.out(wire_94));
  TC_Switch # (.UUID(64'd971606683869478136 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_45 (.en(wire_46), .in(wire_19[15:0]), .out(wire_15_12));
  TC_Switch # (.UUID(64'd488700789590138722 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_46 (.en(wire_73), .in(wire_59[15:0]), .out(wire_24_12));
  TC_Constant # (.UUID(64'd1219804294531623130 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h0)) Constant16_47 (.out(wire_14));
  TC_Switch # (.UUID(64'd2854432665896608476 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_48 (.en(wire_103), .in(wire_127), .out(wire_121));
  TC_Not # (.UUID(64'd1919204710248089503 ^ UUID), .BIT_WIDTH(64'd1)) Not_49 (.in(wire_12), .out(wire_103));
  TC_Switch # (.UUID(64'd3648642341737646920 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_50 (.en(wire_8), .in(wire_2[15:0]), .out(wire_63));
  TC_Switch # (.UUID(64'd2839537485959427856 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_51 (.en(wire_0), .in(wire_0), .out(wire_8));
  TC_Splitter16 # (.UUID(64'd4451072885120255536 ^ UUID)) Splitter16_52 (.in(wire_18[15:0]), .out0(wire_124), .out1());
  TC_Splitter8 # (.UUID(64'd1191888651688547656 ^ UUID)) Splitter8_53 (.in(wire_124), .out0(wire_120), .out1(wire_89), .out2(wire_123), .out3(wire_115), .out4(), .out5(), .out6(), .out7());
  TC_Not # (.UUID(64'd4189336834672528069 ^ UUID), .BIT_WIDTH(64'd1)) Not_54 (.in(wire_6), .out(wire_3));
  TC_Add # (.UUID(64'd3182557287143411779 ^ UUID), .BIT_WIDTH(64'd16)) Add16_55 (.in0(wire_24), .in1(wire_15), .ci(1'd0), .out(wire_33), .co());
  TC_Add # (.UUID(64'd1424675120960351269 ^ UUID), .BIT_WIDTH(64'd16)) Add16_56 (.in0(wire_24), .in1(wire_2[15:0]), .ci(1'd0), .out(wire_77), .co());
  TC_Switch # (.UUID(64'd284020542177892273 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_57 (.en(wire_57), .in(wire_33), .out(wire_1_0));
  TC_Switch # (.UUID(64'd1034703434088870431 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_58 (.en(wire_62), .in(wire_77), .out(wire_1_1));
  TC_Or # (.UUID(64'd657814780105628035 ^ UUID), .BIT_WIDTH(64'd1)) Or_59 (.in0(wire_0), .in1(wire_62), .out(wire_49));
  TC_Console # (.UUID(64'd1550364046122691923 ^ UUID)) Console_60 (.clk(clk), .rst(rst), .offset({{16{1'b0}}, wire_78 }));
  DEC4 # (.UUID(64'd606098422439323267 ^ UUID)) DEC4_61 (.clk(clk), .rst(rst), .Bit_1(wire_111), .Bit_2(wire_118), .Bit_3(wire_67), .Bit_4(wire_128), .Disable(wire_73), .Output_1(wire_5), .Output_2(wire_47), .Output_3(wire_4), .Output_4(wire_23), .Output_5(wire_55), .Output_6(wire_88), .Output_7(wire_97), .Output_8(wire_64), .Output_9(wire_83), .Output_10(wire_65), .Output_11(wire_32), .Output_12(wire_37), .Output_13(), .Output_14(), .Output_15(), .Output_16());
  DEC4 # (.UUID(64'd2350125178974466839 ^ UUID)) DEC4_62 (.clk(clk), .rst(rst), .Bit_1(wire_60), .Bit_2(wire_114), .Bit_3(wire_79), .Bit_4(wire_71), .Disable(wire_46), .Output_1(wire_53), .Output_2(wire_69), .Output_3(wire_51), .Output_4(wire_22), .Output_5(wire_9), .Output_6(wire_11), .Output_7(wire_80), .Output_8(wire_43), .Output_9(wire_29), .Output_10(wire_48), .Output_11(wire_66), .Output_12(wire_40), .Output_13(), .Output_14(), .Output_15(), .Output_16());
  DEC4 # (.UUID(64'd4239434022177334522 ^ UUID)) DEC4_63 (.clk(clk), .rst(rst), .Bit_1(wire_93), .Bit_2(wire_119), .Bit_3(wire_104), .Bit_4(wire_112), .Disable(wire_49), .Output_1(wire_58), .Output_2(wire_42), .Output_3(wire_38), .Output_4(wire_20), .Output_5(wire_16), .Output_6(wire_41), .Output_7(wire_56), .Output_8(wire_61), .Output_9(wire_52), .Output_10(wire_36), .Output_11(wire_26), .Output_12(wire_82), .Output_13(), .Output_14(), .Output_15(), .Output_16());
  DEC2 # (.UUID(64'd2289023201248810830 ^ UUID)) DEC2_64 (.clk(clk), .rst(rst), .Input_1(wire_125), .Input_2(wire_44), .Disable(wire_12), .Output_1(wire_101), .Output_2(wire_6), .Output_3(wire_34), .Output_4(wire_45));
  DEC4 # (.UUID(64'd2197146422829533631 ^ UUID)) DEC4_65 (.clk(clk), .rst(rst), .Bit_1(wire_120), .Bit_2(wire_89), .Bit_3(wire_123), .Bit_4(wire_115), .Disable(wire_3), .Output_1(), .Output_2(), .Output_3(), .Output_4(), .Output_5(), .Output_6(), .Output_7(wire_62), .Output_8(wire_57), .Output_9(), .Output_10(), .Output_11(), .Output_12(), .Output_13(), .Output_14(), .Output_15(), .Output_16());
  ALU # (.UUID(64'd2893949216972807263 ^ UUID)) ALU_66 (.clk(clk), .rst(rst), .Instruction(wire_18[15:0]), .Input_1(wire_24), .Input_2(wire_15), .Enable(wire_45), .Output(wire_30_0[15:0]));
  COND # (.UUID(64'd1476889620975298455 ^ UUID)) COND_67 (.clk(clk), .rst(rst), .Instruction(wire_18[15:0]), .Input_1(wire_24), .Input_2(wire_15), .Enable(wire_101), .Output(wire_0));
  TC_Ram # (.UUID(64'd2067412014399195219 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd65536)) Ram_68 (.clk(clk), .rst(rst), .load(1'd0), .save(wire_39), .address({{16{1'b0}}, wire_24 }), .in0({{48{1'b0}}, wire_15 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(), .out1(), .out2(), .out3());
  TC_Ram # (.UUID(64'd2804227458846121453 ^ UUID), .WORD_WIDTH(64'd16), .WORD_COUNT(64'd32768)) Ram_69 (.clk(clk), .rst(rst), .load(wire_129), .save(wire_1[0:0]), .address({{16{1'b0}}, wire_15 }), .in0(64'd0), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(), .out1(), .out2(), .out3());
  TC_Splitter16 # (.UUID(64'd763171029710359662 ^ UUID)) Splitter16_70 (.in(wire_1), .out0(), .out1(wire_116));
  TC_Splitter8 # (.UUID(64'd3824024877144842064 ^ UUID)) Splitter8_71 (.in(wire_116), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7(wire_28));
  TC_Decoder1 # (.UUID(64'd4576965811034017994 ^ UUID)) Decoder1_72 (.sel(wire_28), .out0(wire_100), .out1(wire_54));
  TC_Switch # (.UUID(64'd2746301141431459897 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_73 (.en(wire_100), .in(wire_62), .out(wire_113));
  TC_Switch # (.UUID(64'd3430101359472696647 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_74 (.en(wire_100), .in(wire_57), .out(wire_81));
  TC_Switch # (.UUID(64'd1728891745001622010 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_75 (.en(wire_54), .in(wire_57), .out(wire_7));
  TC_Switch # (.UUID(64'd4375680025586519226 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_76 (.en(wire_54), .in(wire_62), .out(wire_129));
  TC_Register # (.UUID(64'd2693553474459199961 ^ UUID), .BIT_WIDTH(64'd16)) Register16_77 (.clk(clk), .rst(rst), .load(wire_122), .save(wire_75), .in(wire_85), .out(wire_78));
  TC_Add # (.UUID(64'd3809269893433252203 ^ UUID), .BIT_WIDTH(64'd16)) Add16_78 (.in0(wire_78), .in1(wire_96), .ci(1'd0), .out(wire_85), .co());
  TC_Constant # (.UUID(64'd2151188605745524424 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_79 (.out(wire_122));
  TC_Constant # (.UUID(64'd1918094738540249611 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h50)) Constant16_80 (.out(wire_96));
  TC_Splitter16 # (.UUID(64'd4494426812884145071 ^ UUID)) Splitter16_81 (.in(wire_18[15:0]), .out0(wire_106), .out1());
  TC_Splitter8 # (.UUID(64'd1684985711211094078 ^ UUID)) Splitter8_82 (.in(wire_106), .out0(wire_84), .out1(wire_95), .out2(wire_31), .out3(wire_91), .out4(), .out5(), .out6(), .out7());
  TC_Not # (.UUID(64'd2891551810552540629 ^ UUID), .BIT_WIDTH(64'd1)) Not_83 (.in(wire_34), .out(wire_130));
  DEC4 # (.UUID(64'd2773479126471196673 ^ UUID)) DEC4_84 (.clk(clk), .rst(rst), .Bit_1(wire_84), .Bit_2(wire_95), .Bit_3(wire_31), .Bit_4(wire_91), .Disable(wire_130), .Output_1(), .Output_2(), .Output_3(), .Output_4(), .Output_5(), .Output_6(), .Output_7(wire_75), .Output_8(wire_39), .Output_9(), .Output_10(), .Output_11(), .Output_12(), .Output_13(), .Output_14(), .Output_15(), .Output_16());
  TC_Register # (.UUID(64'd3266843945445956355 ^ UUID), .BIT_WIDTH(64'd16)) Register16_85 (.clk(clk), .rst(rst), .load(wire_70), .save(wire_52), .in(wire_30[15:0]), .out(wire_10));
  TC_Register # (.UUID(64'd373441705232759894 ^ UUID), .BIT_WIDTH(64'd16)) Register16_86 (.clk(clk), .rst(rst), .load(wire_25), .save(wire_36), .in(wire_30[15:0]), .out(wire_72));
  TC_Register # (.UUID(64'd898762616312898673 ^ UUID), .BIT_WIDTH(64'd16)) Register16_87 (.clk(clk), .rst(rst), .load(wire_102), .save(wire_26), .in(wire_30[15:0]), .out(wire_90));
  TC_Register # (.UUID(64'd35259159018310512 ^ UUID), .BIT_WIDTH(64'd16)) Register16_88 (.clk(clk), .rst(rst), .load(wire_74), .save(wire_82), .in(wire_30[15:0]), .out(wire_108));
  TC_Or # (.UUID(64'd3408749404784824565 ^ UUID), .BIT_WIDTH(64'd1)) Or_89 (.in0(wire_83), .in1(wire_29), .out(wire_70));
  TC_Or # (.UUID(64'd2045434085000650231 ^ UUID), .BIT_WIDTH(64'd1)) Or_90 (.in0(wire_65), .in1(wire_48), .out(wire_25));
  TC_Or # (.UUID(64'd4235778316917593708 ^ UUID), .BIT_WIDTH(64'd1)) Or_91 (.in0(wire_32), .in1(wire_66), .out(wire_102));
  TC_Or # (.UUID(64'd1881922342948910945 ^ UUID), .BIT_WIDTH(64'd1)) Or_92 (.in0(wire_37), .in1(wire_40), .out(wire_74));
  TC_Switch # (.UUID(64'd3154836780073834162 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_93 (.en(wire_29), .in(wire_10), .out(wire_15_0));
  TC_Switch # (.UUID(64'd3206739131565530044 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_94 (.en(wire_83), .in(wire_10), .out(wire_24_3));
  TC_Switch # (.UUID(64'd1476550871400967823 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_95 (.en(wire_48), .in(wire_72), .out(wire_15_2));
  TC_Switch # (.UUID(64'd1622071797847061869 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_96 (.en(wire_65), .in(wire_72), .out(wire_24_2));
  TC_Switch # (.UUID(64'd189967047438908968 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_97 (.en(wire_66), .in(wire_90), .out(wire_15_4));
  TC_Switch # (.UUID(64'd3142169352616083849 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_98 (.en(wire_32), .in(wire_90), .out(wire_24_1));
  TC_Switch # (.UUID(64'd2790449206563351533 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_99 (.en(wire_40), .in(wire_108), .out(wire_15_6));
  TC_Switch # (.UUID(64'd1382504743536358321 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_100 (.en(wire_37), .in(wire_108), .out(wire_24_0));

  wire [0:0] wire_0;
  wire [15:0] wire_1;
  wire [15:0] wire_1_0;
  wire [15:0] wire_1_1;
  assign wire_1 = wire_1_0|wire_1_1;
  wire [63:0] wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [15:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [7:0] wire_13;
  wire [15:0] wire_14;
  wire [15:0] wire_15;
  wire [15:0] wire_15_0;
  wire [15:0] wire_15_1;
  wire [15:0] wire_15_2;
  wire [15:0] wire_15_3;
  wire [15:0] wire_15_4;
  wire [15:0] wire_15_5;
  wire [15:0] wire_15_6;
  wire [15:0] wire_15_7;
  wire [15:0] wire_15_8;
  wire [15:0] wire_15_9;
  wire [15:0] wire_15_10;
  wire [15:0] wire_15_11;
  wire [15:0] wire_15_12;
  assign wire_15 = wire_15_0|wire_15_1|wire_15_2|wire_15_3|wire_15_4|wire_15_5|wire_15_6|wire_15_7|wire_15_8|wire_15_9|wire_15_10|wire_15_11|wire_15_12;
  wire [0:0] wire_16;
  wire [15:0] wire_17;
  wire [63:0] wire_18;
  wire [63:0] wire_19;
  wire [0:0] wire_20;
  wire [15:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [15:0] wire_24;
  wire [15:0] wire_24_0;
  wire [15:0] wire_24_1;
  wire [15:0] wire_24_2;
  wire [15:0] wire_24_3;
  wire [15:0] wire_24_4;
  wire [15:0] wire_24_5;
  wire [15:0] wire_24_6;
  wire [15:0] wire_24_7;
  wire [15:0] wire_24_8;
  wire [15:0] wire_24_9;
  wire [15:0] wire_24_10;
  wire [15:0] wire_24_11;
  wire [15:0] wire_24_12;
  assign wire_24 = wire_24_0|wire_24_1|wire_24_2|wire_24_3|wire_24_4|wire_24_5|wire_24_6|wire_24_7|wire_24_8|wire_24_9|wire_24_10|wire_24_11|wire_24_12;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [63:0] wire_30;
  wire [63:0] wire_30_0;
  wire [63:0] wire_30_1;
  assign wire_30 = wire_30_0|wire_30_1;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [15:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [0:0] wire_58;
  wire [63:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [15:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [15:0] wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [15:0] wire_72;
  wire [0:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [15:0] wire_76;
  wire [15:0] wire_77;
  wire [15:0] wire_78;
  wire [0:0] wire_79;
  wire [0:0] wire_80;
  wire [0:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;
  wire [0:0] wire_84;
  wire [15:0] wire_85;
  wire [15:0] wire_86;
  wire [7:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;
  wire [15:0] wire_90;
  wire [0:0] wire_91;
  wire [0:0] wire_92;
  wire [0:0] wire_93;
  wire [15:0] wire_94;
  wire [0:0] wire_95;
  wire [15:0] wire_96;
  wire [0:0] wire_97;
  wire [15:0] wire_98;
  wire [0:0] wire_99;
  wire [0:0] wire_100;
  wire [0:0] wire_101;
  wire [0:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [0:0] wire_105;
  wire [7:0] wire_106;
  wire [0:0] wire_107;
  wire [15:0] wire_108;
  wire [7:0] wire_109;
  wire [0:0] wire_110;
  wire [0:0] wire_111;
  wire [0:0] wire_112;
  wire [0:0] wire_113;
  wire [0:0] wire_114;
  wire [0:0] wire_115;
  wire [7:0] wire_116;
  wire [15:0] wire_117;
  wire [0:0] wire_118;
  wire [0:0] wire_119;
  wire [0:0] wire_120;
  wire [7:0] wire_121;
  wire [0:0] wire_122;
  wire [0:0] wire_123;
  wire [7:0] wire_124;
  wire [0:0] wire_125;
  wire [15:0] wire_126;
  wire [7:0] wire_127;
  wire [0:0] wire_128;
  wire [0:0] wire_129;
  wire [0:0] wire_130;

endmodule
