module ALU (clk, rst, Instruction, Input_1, Input_2, Enable, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [15:0] Instruction;
  input  wire [15:0] Input_1;
  input  wire [15:0] Input_2;
  input  wire [0:0] Enable;
  output  wire [15:0] Output;

  TC_Splitter16 # (.UUID(64'd129274797608114045 ^ UUID)) Splitter16_0 (.in(wire_9), .out0(wire_14), .out1());
  TC_Splitter8 # (.UUID(64'd1462455766308944097 ^ UUID)) Splitter8_1 (.in(wire_14), .out0(wire_20), .out1(wire_5), .out2(wire_34), .out3(wire_37), .out4(), .out5(), .out6(), .out7());
  TC_Add # (.UUID(64'd960219409565390549 ^ UUID), .BIT_WIDTH(64'd16)) Add16_2 (.in0(wire_11), .in1(wire_2), .ci(1'd0), .out(wire_38), .co());
  TC_Add # (.UUID(64'd3710995179557622515 ^ UUID), .BIT_WIDTH(64'd16)) Add16_3 (.in0(wire_11), .in1(wire_35), .ci(1'd0), .out(wire_19), .co());
  TC_Mul # (.UUID(64'd2979747764176318793 ^ UUID), .BIT_WIDTH(64'd16)) Mul16_4 (.in0(wire_11), .in1(wire_2), .out0(wire_29), .out1());
  TC_Mul # (.UUID(64'd4112779538525025640 ^ UUID), .BIT_WIDTH(64'd16)) DivMod16_5 (.in0(wire_11), .in1(wire_1), .out0(wire_33), .out1(wire_27));
  TC_Neg # (.UUID(64'd2530762749794426659 ^ UUID), .BIT_WIDTH(64'd16)) Neg16_6 (.in(wire_2), .out(wire_35));
  TC_Shl # (.UUID(64'd3696538209267226338 ^ UUID), .BIT_WIDTH(64'd16)) Shl16_7 (.in(wire_11), .shift(wire_2[7:0]), .out(wire_0));
  TC_Shr # (.UUID(64'd558338407377449065 ^ UUID), .BIT_WIDTH(64'd16)) Shr16_8 (.in(wire_11), .shift(wire_2[7:0]), .out(wire_25));
  TC_Ashr # (.UUID(64'd749026858371219188 ^ UUID), .BIT_WIDTH(64'd16)) Ashr16_9 (.in(wire_11), .shift(wire_2[7:0]), .out(wire_36));
  TC_And # (.UUID(64'd3902266159717928988 ^ UUID), .BIT_WIDTH(64'd16)) And16_10 (.in0(wire_11), .in1(wire_2), .out(wire_32));
  TC_Or # (.UUID(64'd1626630594968710822 ^ UUID), .BIT_WIDTH(64'd16)) Or16_11 (.in0(wire_11), .in1(wire_2), .out(wire_22));
  TC_Xor # (.UUID(64'd108456683173740732 ^ UUID), .BIT_WIDTH(64'd16)) Xor16_12 (.in0(wire_11), .in1(wire_2), .out(wire_17));
  TC_Not # (.UUID(64'd1072175468325980639 ^ UUID), .BIT_WIDTH(64'd16)) Not16_13 (.in(wire_11), .out(wire_4));
  TC_Switch # (.UUID(64'd1106245126962629211 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_14 (.en(wire_28), .in(wire_38), .out(wire_6_3));
  TC_Switch # (.UUID(64'd1699455517898077188 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_15 (.en(wire_30), .in(wire_19), .out(wire_6_2));
  TC_Switch # (.UUID(64'd1037848991120861857 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_16 (.en(wire_16), .in(wire_29), .out(wire_6_0));
  TC_Switch # (.UUID(64'd2679548854247736178 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_17 (.en(wire_10), .in(wire_33), .out(wire_6_1));
  TC_Switch # (.UUID(64'd664042728090713532 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_18 (.en(wire_23), .in(wire_0), .out(wire_6_5));
  TC_Switch # (.UUID(64'd1773019090982858830 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_19 (.en(wire_31), .in(wire_25), .out(wire_6_6));
  TC_Switch # (.UUID(64'd1527054064579548263 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_20 (.en(wire_21), .in(wire_27), .out(wire_6_4));
  TC_Switch # (.UUID(64'd3230975643929287438 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_21 (.en(wire_13), .in(wire_36), .out(wire_6_7));
  TC_Switch # (.UUID(64'd2364361064743946803 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_22 (.en(wire_24), .in(wire_32), .out(wire_6_8));
  TC_Switch # (.UUID(64'd3178299767776664427 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_23 (.en(wire_3), .in(wire_22), .out(wire_6_9));
  TC_Switch # (.UUID(64'd2635356813930944275 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_24 (.en(wire_18), .in(wire_17), .out(wire_6_10));
  TC_Switch # (.UUID(64'd2650181991435326595 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_25 (.en(wire_15), .in(wire_4), .out(wire_6_11));
  TC_Maker16 # (.UUID(64'd4157917437721305216 ^ UUID)) Maker16_26 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd2530465127559157045 ^ UUID)) Maker16_27 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd3318448313327833152 ^ UUID)) Maker16_28 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd1341563485140346365 ^ UUID)) Maker16_29 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd2448306895543285647 ^ UUID)) Maker16_30 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd2982555009944348411 ^ UUID)) Maker16_31 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd3715244167020249352 ^ UUID)) Maker16_32 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd795844953056343003 ^ UUID)) Maker16_33 (.in0(8'd0), .in1(8'd0), .out());
  TC_Not # (.UUID(64'd1276716563455362769 ^ UUID), .BIT_WIDTH(64'd1)) Not_34 (.in(1'd0), .out());
  TC_Not # (.UUID(64'd3642479983096000307 ^ UUID), .BIT_WIDTH(64'd1)) Not_35 (.in(1'd0), .out());
  TC_Switch # (.UUID(64'd557744667485185326 ^ UUID), .BIT_WIDTH(64'd16)) Output16z_36 (.en(wire_26), .in(wire_6), .out(Output));
  TC_Equal # (.UUID(64'd2494304255186729504 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_37 (.in0(wire_2), .in1(16'd0), .out(wire_8));
  TC_Not # (.UUID(64'd2360878654635395758 ^ UUID), .BIT_WIDTH(64'd1)) Not_38 (.in(wire_8), .out(wire_7));
  TC_Switch # (.UUID(64'd47150918006556051 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_39 (.en(wire_8), .in(wire_12), .out(wire_1_1));
  TC_Constant # (.UUID(64'd3324600182956937994 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h1)) Constant16_40 (.out(wire_12));
  TC_Switch # (.UUID(64'd3951192607140037191 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_41 (.en(wire_7), .in(wire_2), .out(wire_1_0));
  DEC4 # (.UUID(64'd1718291227987089359 ^ UUID)) DEC4_42 (.clk(clk), .rst(rst), .Bit_1(wire_20), .Bit_2(wire_5), .Bit_3(wire_34), .Bit_4(wire_37), .Disable(1'd0), .Output_1(wire_23), .Output_2(wire_31), .Output_3(wire_13), .Output_4(wire_21), .Output_5(wire_10), .Output_6(wire_16), .Output_7(wire_30), .Output_8(wire_28), .Output_9(wire_24), .Output_10(wire_3), .Output_11(wire_18), .Output_12(wire_15), .Output_13(), .Output_14(), .Output_15(), .Output_16());

  wire [15:0] wire_0;
  wire [15:0] wire_1;
  wire [15:0] wire_1_0;
  wire [15:0] wire_1_1;
  assign wire_1 = wire_1_0|wire_1_1;
  wire [15:0] wire_2;
  assign wire_2 = Input_2;
  wire [0:0] wire_3;
  wire [15:0] wire_4;
  wire [0:0] wire_5;
  wire [15:0] wire_6;
  wire [15:0] wire_6_0;
  wire [15:0] wire_6_1;
  wire [15:0] wire_6_2;
  wire [15:0] wire_6_3;
  wire [15:0] wire_6_4;
  wire [15:0] wire_6_5;
  wire [15:0] wire_6_6;
  wire [15:0] wire_6_7;
  wire [15:0] wire_6_8;
  wire [15:0] wire_6_9;
  wire [15:0] wire_6_10;
  wire [15:0] wire_6_11;
  assign wire_6 = wire_6_0|wire_6_1|wire_6_2|wire_6_3|wire_6_4|wire_6_5|wire_6_6|wire_6_7|wire_6_8|wire_6_9|wire_6_10|wire_6_11;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [15:0] wire_9;
  assign wire_9 = Instruction;
  wire [0:0] wire_10;
  wire [15:0] wire_11;
  assign wire_11 = Input_1;
  wire [15:0] wire_12;
  wire [0:0] wire_13;
  wire [7:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [15:0] wire_17;
  wire [0:0] wire_18;
  wire [15:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [15:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [15:0] wire_25;
  wire [0:0] wire_26;
  assign wire_26 = Enable;
  wire [15:0] wire_27;
  wire [0:0] wire_28;
  wire [15:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [15:0] wire_32;
  wire [15:0] wire_33;
  wire [0:0] wire_34;
  wire [15:0] wire_35;
  wire [15:0] wire_36;
  wire [0:0] wire_37;
  wire [15:0] wire_38;

endmodule
