module OPP8 (clk, rst, Input_1, Input_2, Input_3, Input_4, Input_5, Input_6, Input_7, Input_8, Enable_All, Output_1, Output_2, Output_3, Output_4, Output_5, Output_6, Output_7, Output_8);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] Input_1;
  input  wire [0:0] Input_2;
  input  wire [0:0] Input_3;
  input  wire [0:0] Input_4;
  input  wire [0:0] Input_5;
  input  wire [0:0] Input_6;
  input  wire [0:0] Input_7;
  input  wire [0:0] Input_8;
  input  wire [0:0] Enable_All;
  output  wire [0:0] Output_1;
  output  wire [0:0] Output_2;
  output  wire [0:0] Output_3;
  output  wire [0:0] Output_4;
  output  wire [0:0] Output_5;
  output  wire [0:0] Output_6;
  output  wire [0:0] Output_7;
  output  wire [0:0] Output_8;

  TC_Maker16 # (.UUID(64'd4576894713119714030 ^ UUID)) Maker16_0 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd4159457257671284809 ^ UUID)) Maker16_1 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd135754618811469109 ^ UUID)) Maker16_2 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd2144888840407442937 ^ UUID)) Maker16_3 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd1923742623033063111 ^ UUID)) Maker16_4 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd2531585302615411283 ^ UUID)) Maker16_5 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd1446271324425451477 ^ UUID)) Maker16_6 (.in0(8'd0), .in1(8'd0), .out());
  TC_Maker16 # (.UUID(64'd971499438910037494 ^ UUID)) Maker16_7 (.in0(8'd0), .in1(8'd0), .out());
  TC_Or # (.UUID(64'd2495172288979506291 ^ UUID), .BIT_WIDTH(64'd1)) Or_8 (.in0(wire_1), .in1(wire_5), .out(wire_10));
  TC_Or # (.UUID(64'd501113617363284001 ^ UUID), .BIT_WIDTH(64'd1)) Or_9 (.in0(wire_1), .in1(wire_4), .out(wire_12));
  TC_Or # (.UUID(64'd3512947802125280731 ^ UUID), .BIT_WIDTH(64'd1)) Or_10 (.in0(wire_1), .in1(wire_6), .out(wire_15));
  TC_Or # (.UUID(64'd142855482572645156 ^ UUID), .BIT_WIDTH(64'd1)) Or_11 (.in0(wire_1), .in1(wire_9), .out(wire_3));
  TC_Or # (.UUID(64'd1751663132027682070 ^ UUID), .BIT_WIDTH(64'd1)) Or_12 (.in0(wire_1), .in1(wire_7), .out(wire_16));
  TC_Or # (.UUID(64'd3398456072975241789 ^ UUID), .BIT_WIDTH(64'd1)) Or_13 (.in0(wire_1), .in1(wire_2), .out(wire_13));
  TC_Or # (.UUID(64'd885462322106012501 ^ UUID), .BIT_WIDTH(64'd1)) Or_14 (.in0(wire_1), .in1(wire_0), .out(wire_14));
  TC_Or # (.UUID(64'd2601404253331207743 ^ UUID), .BIT_WIDTH(64'd1)) Or_15 (.in0(wire_1), .in1(wire_8), .out(wire_11));

  wire [0:0] wire_0;
  assign wire_0 = Input_2;
  wire [0:0] wire_1;
  assign wire_1 = Enable_All;
  wire [0:0] wire_2;
  assign wire_2 = Input_3;
  wire [0:0] wire_3;
  assign Output_4 = wire_3;
  wire [0:0] wire_4;
  assign wire_4 = Input_7;
  wire [0:0] wire_5;
  assign wire_5 = Input_8;
  wire [0:0] wire_6;
  assign wire_6 = Input_6;
  wire [0:0] wire_7;
  assign wire_7 = Input_4;
  wire [0:0] wire_8;
  assign wire_8 = Input_1;
  wire [0:0] wire_9;
  assign wire_9 = Input_5;
  wire [0:0] wire_10;
  assign Output_1 = wire_10;
  wire [0:0] wire_11;
  assign Output_8 = wire_11;
  wire [0:0] wire_12;
  assign Output_2 = wire_12;
  wire [0:0] wire_13;
  assign Output_6 = wire_13;
  wire [0:0] wire_14;
  assign Output_7 = wire_14;
  wire [0:0] wire_15;
  assign Output_3 = wire_15;
  wire [0:0] wire_16;
  assign Output_5 = wire_16;

endmodule
